module crab (
    input [9:0] h_cnt,
    input [9:0] v_cnt,
    input [9:0] fish_h_position,
    input [9:0] fish_v_position,
    input fish_way,  //0 for go left , 1 for go right
    input appear,
    input type,
    output reg background, //1 for print background 0 for print fish
    output reg [11:0] vga
);
    parameter [11:0] crab1 [0:899] = {//30*30
        //get rid of 353,351,452,453, 463, 464 etc.
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h231,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h252,12'h352,12'h352,12'hE87,12'h621,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h531,12'h441,12'h352,12'hE64,12'hF53,12'h320,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h420,12'hF52,12'hE54,12'h610,12'hF63,12'hF53,12'h931,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h932,12'hF53,12'hF52,12'hF53,12'hF53,12'hF63,12'hC21,12'h341,12'h352,12'h352,
        12'h352,12'h352,12'hB98,12'h352,12'h352,12'h331,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'hB52,12'hE63,12'hF53,12'hF53,12'hF53,12'hF63,12'hD30,12'h330,12'h352,12'h352,
        12'h352,12'h632,12'hF76,12'h341,12'h431,12'hD54,12'h942,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h932,12'hF52,12'hF53,12'hF53,12'hF53,12'hF53,12'hD20,12'h330,12'h352,12'h352,
        12'h352,12'hF54,12'hF53,12'hC65,12'hC53,12'hF53,12'hF53,12'h430,12'h352,12'h352,12'h352,12'h242,12'h352,12'h352,12'h352,12'h352,12'h010,12'h120,12'h352,12'h352,12'h320,12'hF53,12'hF53,12'hF53,12'hF53,12'hE52,12'hC31,12'h341,12'h352,12'h352,
        12'h352,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'h942,12'h352,12'h352,12'h120,12'h120,12'h352,12'h352,12'h352,12'h352,12'h352,12'h341,12'h352,12'h352,12'h352,12'hC43,12'hE42,12'hD31,12'hF53,12'hD30,12'h831,12'h352,12'h352,12'h352,
        12'h352,12'hE42,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hD64,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'hABB,12'h100,12'h565,12'h352,12'h251,12'h431,12'hC32,12'hB30,12'hD20,12'h821,12'h352,12'h352,12'h352,12'h352,
        12'h341,12'hD42,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hE64,12'h242,12'h352,12'h352,12'h010,12'h352,12'h352,12'h352,12'h352,12'hFFF,12'hFFF,12'hEDD,12'h242,12'h252,12'h352,12'h842,12'h400,12'h331,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'hB32,12'hF52,12'hF53,12'hF53,12'hF53,12'hF53,12'h942,12'h352,12'h352,12'h888,12'h889,12'hFFF,12'h865,12'hF87,12'hF66,12'hDCC,12'hFFF,12'h855,12'hE53,12'hF54,12'h721,12'hD53,12'h330,12'h352,12'h341,12'hD53,12'h731,12'h352,12'h352,
        12'h352,12'h410,12'hC31,12'hE41,12'hF53,12'hE53,12'hF53,12'h320,12'h352,12'h352,12'h777,12'hFFF,12'hFFF,12'hD55,12'hF53,12'hF53,12'hD54,12'hB42,12'hF53,12'hF53,12'hF53,12'hF53,12'hC52,12'h352,12'h330,12'hF64,12'hA42,12'hE53,12'h441,12'h352,
        12'h352,12'h352,12'h720,12'hC31,12'hC30,12'hC30,12'h710,12'h352,12'h341,12'hC64,12'hE64,12'h754,12'h621,12'hF63,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'h932,12'hE43,12'hB42,12'h352,12'h320,12'h531,12'h352,
        12'h352,12'h352,12'h352,12'h441,12'h330,12'h410,12'hB53,12'h421,12'hE63,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF63,12'h620,12'h331,12'h352,12'h352,12'h231,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h821,12'hE63,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF42,12'hC43,12'h352,12'h251,12'h331,12'h331,12'h352,
        12'h352,12'h352,12'h442,12'h231,12'h352,12'h352,12'hB53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hE52,12'hD32,12'h932,12'hD42,12'hE63,12'hE53,12'h352,
        12'h352,12'h352,12'h541,12'hF54,12'hA43,12'h331,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF63,12'hE64,12'hF63,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hE52,12'hC21,12'h320,12'h410,12'hA32,12'hE53,12'h441,
        12'h352,12'h352,12'hD53,12'hE63,12'hE32,12'h931,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hE53,12'hE64,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hD31,12'hB31,12'h352,12'h352,12'h352,12'h742,12'h441,
        12'h352,12'h352,12'hC53,12'h352,12'h331,12'h410,12'hF42,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hE53,12'hE54,12'hE64,12'hA21,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hC31,12'hD31,12'h420,12'h352,12'h352,12'h352,12'h432,12'h442,
        12'h352,12'h331,12'h230,12'h352,12'h352,12'h352,12'hD43,12'hF52,12'hF53,12'hF53,12'hF53,12'hF53,12'hE53,12'hE54,12'hE64,12'hB42,12'hD53,12'hF53,12'hF53,12'hF53,12'hF53,12'hE31,12'hC21,12'h600,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h220,12'h352,12'h352,12'h320,12'hC54,12'h820,12'hE41,12'hF52,12'hF53,12'hF53,12'hF53,12'hF64,12'hF64,12'hF53,12'hF52,12'hF53,12'hF53,12'hF53,12'hF52,12'hC30,12'h931,12'h410,12'hD31,12'hA53,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h240,12'h352,12'h421,12'hE63,12'hD31,12'h510,12'hC31,12'hE42,12'hF43,12'hE53,12'hF53,12'hF53,12'hF53,12'hF52,12'hF53,12'hF53,12'hF52,12'hD41,12'hC30,12'h731,12'h331,12'h352,12'h821,12'hE53,12'h510,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h320,12'hF53,12'hE42,12'h320,12'h352,12'h410,12'hC31,12'hC31,12'hC30,12'hD42,12'hE42,12'hE42,12'hE41,12'hD31,12'hC20,12'hB31,12'h520,12'h331,12'h352,12'h352,12'h352,12'h352,12'hF63,12'h520,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h321,12'hF53,12'h310,12'h352,12'h352,12'h331,12'hB43,12'h510,12'hA21,12'hB31,12'hB31,12'h920,12'h410,12'h320,12'h341,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h420,12'h742,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'hF54,12'h341,12'h352,12'h352,12'h731,12'hE41,12'h320,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h421,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'hA53,12'h241,12'h352,12'h352,12'hC53,12'hC42,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h320,12'h332,12'h352,12'h352,12'h420,12'hE64,12'h320,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h361,12'h352,12'h231,12'h352,12'h352,12'h352,12'h431,12'hB54,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h120,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352
    };

    parameter [11:0] crab2 [0:899] = {//30*30
        //get rid of 353,351,452,453, 463, 464 etc.
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h341,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h330,12'hD75,12'h221,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h341,12'hE64,12'hE53,12'h331,12'h352,12'h331,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h720,12'hF53,12'hF53,12'hB43,12'hA42,12'hF54,12'h630,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'hC41,12'hF53,12'hF53,12'hF63,12'hF53,12'hF53,12'hC53,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h241,12'hD42,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hD63,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h231,12'hD31,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hC53,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h341,12'h420,12'h252,12'h352,12'h976,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'hB31,12'hF53,12'hF53,12'hF53,12'hF63,12'hF53,12'h631,12'h352,12'h352,12'h010,12'h231,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'hE53,12'hE53,12'h331,12'h431,12'hE54,12'h430,
        12'h352,12'h352,12'h352,12'h352,12'h721,12'hD31,12'hE52,12'hF53,12'hF53,12'hE64,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h120,12'h352,12'h352,12'h352,12'h731,12'hF53,12'hF53,12'hB31,12'hD53,12'hF53,12'h921,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h921,12'hC31,12'hD31,12'hC41,12'h431,12'h352,12'h352,12'h444,12'h110,12'h343,12'h352,12'h352,12'h352,12'h352,12'h231,12'h242,12'h352,12'h352,12'hE63,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hB32,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h320,12'h500,12'h432,12'h352,12'h352,12'h242,12'hFFF,12'h222,12'h676,12'h352,12'h352,12'h352,12'h121,12'h231,12'h352,12'h352,12'h352,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hC21,
        12'h352,12'h352,12'h352,12'h542,12'h341,12'h352,12'h352,12'hD43,12'h331,12'h831,12'hD75,12'hA54,12'hFFF,12'hFFF,12'h865,12'h964,12'h542,12'h343,12'hCBC,12'h555,12'h352,12'h352,12'h352,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF42,12'hA32,
        12'h352,12'h352,12'h330,12'hF53,12'h941,12'h352,12'h352,12'hA31,12'hF53,12'hF53,12'hF53,12'hF53,12'h732,12'h977,12'hD54,12'hF52,12'hF53,12'hA88,12'hFFF,12'hFFF,12'h352,12'h352,12'h352,12'hC41,12'hE42,12'hF53,12'hF53,12'hF53,12'hC30,12'h510,
        12'h252,12'h352,12'hE54,12'hD63,12'hF53,12'h320,12'hB53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF54,12'hF53,12'hF52,12'hF63,12'hF53,12'hB54,12'hEED,12'hB88,12'h843,12'h352,12'h352,12'h510,12'hE42,12'hD31,12'hE42,12'hD41,12'hC31,12'h341,
        12'h352,12'h632,12'h331,12'h352,12'h820,12'h710,12'hF52,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF54,12'hF53,12'hF63,12'hC53,12'h341,12'h933,12'h920,12'hC31,12'hC31,12'hB31,12'h330,12'h352,
        12'h241,12'h352,12'h352,12'h352,12'h352,12'hA43,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF63,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hB43,12'hD41,12'h242,12'h352,12'h341,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h331,12'h320,12'hB43,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'h310,12'h352,12'h352,12'h352,12'h331,12'h352,12'h352,
        12'h352,12'hA53,12'hE53,12'hF53,12'hE42,12'hB31,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF64,12'hF63,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'h631,12'h420,12'hC54,12'hE54,12'hC54,12'h352,12'h352,
        12'h341,12'hF54,12'hE53,12'h620,12'h320,12'h731,12'hE42,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hE64,12'hE54,12'hE54,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF52,12'hD53,12'hD42,12'hB42,12'h310,12'hF63,12'h352,12'h352,
        12'h352,12'hF53,12'h431,12'h352,12'h251,12'h430,12'hC21,12'hE52,12'hF53,12'hF53,12'hE64,12'hE54,12'hE64,12'hB53,12'hF64,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hE53,12'h520,12'h352,12'h352,12'h731,12'h252,12'h352,
        12'h341,12'hD53,12'h352,12'h352,12'h352,12'h320,12'h810,12'hC30,12'hD41,12'hF53,12'hF63,12'hF63,12'hF64,12'hD63,12'hA21,12'hE53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hE42,12'hE43,12'h352,12'h352,12'h252,12'h332,12'h352,12'h352,
        12'h441,12'h310,12'h352,12'h352,12'h441,12'hE53,12'hB32,12'h831,12'hD21,12'hD31,12'hF52,12'hF53,12'hF53,12'hF53,12'hE53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hF53,12'hD31,12'hA30,12'hB42,12'hA42,12'h420,12'h352,12'h352,12'h352,
        12'h341,12'h331,12'h352,12'h352,12'h731,12'hD42,12'h320,12'h241,12'h720,12'hC31,12'hC31,12'hF42,12'hF53,12'hF53,12'hF53,12'hF52,12'hF53,12'hF53,12'hF53,12'hF53,12'hE52,12'hE31,12'hD20,12'h510,12'h921,12'hE41,12'hE53,12'h732,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h832,12'h820,12'h352,12'h352,12'h252,12'h431,12'h510,12'hA31,12'hB21,12'hD30,12'hE42,12'hF53,12'hF53,12'hF53,12'hF53,12'hE32,12'hD20,12'hC31,12'h921,12'h352,12'h352,12'h610,12'hF53,12'h932,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h331,12'hC54,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h341,12'h310,12'h621,12'h931,12'hB31,12'hB31,12'hB31,12'hA31,12'h820,12'h210,12'h352,12'h352,12'h352,12'h352,12'hA33,12'h331,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h621,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'hA32,12'hC53,12'h352,12'h352,12'h352,12'h352,12'h854,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h442,12'h010,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h520,12'hF43,12'h331,12'h352,12'h352,12'h352,12'h341,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h932,12'hE64,12'h331,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h632,12'h520,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352
    };


    always @(*) begin
        background = 1'b1;
        vga = 12'h000;
        if(appear == 1'b0) begin
            background = 1'b1;
            vga = 12'h000;
        end
        else if(type == 1'b0) begin
            if(((h_cnt+30) - fish_h_position) <= 29 && (v_cnt - fish_v_position) <= 29) begin
                if(crab1[(v_cnt - fish_v_position) * 30 + (h_cnt + 30 - fish_h_position)] != 12'h352) begin
                    background = 0;
                    vga = crab1[(v_cnt - fish_v_position) * 30 + (h_cnt + 30 - fish_h_position)];
                end
                else begin
                    background = 1;
                    vga = 12'h000;
                end
            end
            else begin
                background = 1;
                vga = 12'h000;
            end
        end
        else if(type == 1'b1) begin
            if(((h_cnt+30) - fish_h_position) <= 29 && (v_cnt - fish_v_position) <= 29) begin
                if(crab2[(v_cnt - fish_v_position) * 30 + (h_cnt + 30 - fish_h_position)] != 12'h352) begin
                    background = 0;
                    vga = crab2[(v_cnt - fish_v_position) * 30 + (h_cnt + 30 - fish_h_position)];
                end
                else begin
                    background = 1;
                    vga = 12'h000;
                end
            end
            else begin
                background = 1;
                vga = 12'h000;
            end
        end
        else begin
            background = 1;
            vga = 12'h000;
        end


    end
    
endmodule


        