
module play (
    input [9:0] h_cnt,
    input [9:0] v_cnt,
    output reg background, //1 for print background 0 for print fish
    output reg [11:0] vga
);
    parameter [11:0] play [0:2399] = {//60*40
    
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hADF,12'hAEF,12'hAEF,12'hAEF,12'hADF,12'hAEF,12'hAEF,12'hAEF,12'hADF,12'hAEF,12'h9EF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEE,12'hAEF,12'hAEF,12'hADF,12'hADF,12'hADF,12'hAEF,12'hAEF,12'hADF,12'hADF,12'hAEF,12'hAEF,12'hAEE,12'hAEF,12'hAEF,12'hADF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hADF,12'hAEF,12'hAEF,12'hADF,12'hAEF,12'hAEE,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'h9EF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hADF,12'hBDF,12'hBDE,12'hACC,12'hACC,12'hADD,12'hAEE,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'h9EF,12'hAEF,12'hAEF,12'hAEF,12'hBDE,12'hACC,12'hBCC,12'hACC,12'hBDE,12'hAEE,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEE,12'hBDD,12'hAB8,12'hAA6,12'hBC9,12'hCC9,12'hDDA,12'hDB8,12'hA97,12'hAB8,12'hADC,12'hADD,12'hAEE,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hADF,12'hADF,12'hBDE,12'hADC,12'hAA8,12'hAA7,12'hDC9,12'hDD9,12'hCC9,12'hBB8,12'hAA7,12'hBB9,12'hACC,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEE,12'h9BA,12'hBB8,12'hFEC,12'hFFF,12'hFFE,12'hFFE,12'hFFF,12'hFFF,12'hFFE,12'hFFD,12'hDC8,12'hAA7,12'hAB9,12'hACC,12'hADD,12'hADE,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hADF,12'hADD,12'hBCB,12'hAB8,12'hBA7,12'hDC9,12'hFFD,12'hFFE,12'hFFF,12'hFFF,12'hFFF,12'hFFE,12'hFFE,12'hFFC,12'hBB7,12'hBA8,12'hAEE,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAB9,12'hEEB,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFC,12'hFEB,12'hFFC,12'hFFE,12'hFFF,12'hFFF,12'hFFE,12'hFFD,12'hEEB,12'hBB9,12'h997,12'hAB9,12'hABA,12'hBCB,12'hBCC,12'hBDD,12'hAEF,12'hADF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBEE,12'hBDE,12'hBDD,12'hABA,12'hABA,12'hAB9,12'hBB8,12'hEDB,12'hFFD,12'hFFE,12'hFFE,12'hFFE,12'hFFD,12'hFFB,12'hFEB,12'hFFB,12'hFFC,12'hFFE,12'hFFF,12'hFFE,12'hEEB,12'hAA8,12'hAEE,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBCB,12'hEEA,12'hFFF,12'hFFE,12'hEEB,12'hEEB,12'hFFC,12'hED9,12'hEC6,12'hEC5,12'hED6,12'hFD8,12'hFFB,12'hFFD,12'hFFE,12'hFFF,12'hFFE,12'hFFE,12'hFFD,12'hFEB,12'hDC9,12'hCB8,12'hAA7,12'hAA8,12'hAA8,12'hAA7,12'hAA7,12'hAA7,12'hAA8,12'hBA8,12'hCB9,12'hDCA,12'hFEB,12'hFFD,12'hFFE,12'hFFE,12'hFFF,12'hFFE,12'hFFD,12'hFEA,12'hED8,12'hEC6,12'hEC5,12'hEC5,12'hEC5,12'hEC5,12'hEC6,12'hED9,12'hFFC,12'hFFE,12'hFEB,12'hAB9,12'hADF,12'hAEF,12'hAEF,12'hAEF,
        12'hADF,12'hAEF,12'hAEF,12'hADF,12'hAA6,12'hFFF,12'hFFC,12'hDD7,12'hFEB,12'hFFD,12'hFFE,12'hFFE,12'hED7,12'hFC3,12'hFC4,12'hFC5,12'hEC5,12'hEC6,12'hED8,12'hFEA,12'hFFC,12'hFFD,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFE,12'hFFE,12'hFFD,12'hFFD,12'hFFD,12'hFFD,12'hFFE,12'hFFE,12'hFFE,12'hFFF,12'hFFF,12'hFFF,12'hFFD,12'hFFC,12'hFEA,12'hED7,12'hEC6,12'hEC5,12'hEC4,12'hFC4,12'hFC4,12'hFC4,12'hFC4,12'hFD4,12'hFC4,12'hEB2,12'hDB4,12'hFFC,12'hFFE,12'hDC9,12'hADD,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hBDC,12'hFEC,12'hFFE,12'hFD7,12'hED7,12'hFFD,12'hFFE,12'hFFE,12'hFFF,12'hFFA,12'hFD4,12'hFD4,12'hEC4,12'hFC4,12'hFC4,12'hFC5,12'hFC5,12'hEC5,12'hEC6,12'hED8,12'hFD9,12'hFEA,12'hFFC,12'hFFD,12'hFFE,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFE,12'hFFD,12'hFFD,12'hFFB,12'hFE9,12'hED8,12'hED6,12'hEC5,12'hEC5,12'hFC4,12'hFC4,12'hFC4,12'hFC4,12'hEC4,12'hFC4,12'hFD4,12'hFD4,12'hFC4,12'hEC2,12'hEB2,12'hEB2,12'hDB4,12'hFFD,12'hFFE,12'h9A8,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hADF,12'h9A7,12'hFFF,12'hFFB,12'hEC5,12'hFE9,12'hFFE,12'hFFE,12'hFFE,12'hFFD,12'hFE9,12'hFE5,12'hFE5,12'hFE5,12'hFD5,12'hFD4,12'hEC4,12'hEC4,12'hFC4,12'hFC4,12'hEC4,12'hEC4,12'hEC5,12'hEC6,12'hEC6,12'hEC6,12'hEC6,12'hEC6,12'hED7,12'hEC6,12'hEC6,12'hED5,12'hED5,12'hED5,12'hEC5,12'hED4,12'hEC4,12'hEC3,12'hED4,12'hFC5,12'hFC4,12'hFD4,12'hFD5,12'hFE5,12'hFE5,12'hFE4,12'hFD4,12'hFD4,12'hFD4,12'hEC2,12'hEB2,12'hEB2,12'hDC6,12'hFFF,12'hCB8,12'hAEE,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hADF,12'hAB7,12'hFFE,12'hFE8,12'hEC5,12'hFEA,12'hFFE,12'hFFE,12'hFFD,12'hFFA,12'hFE6,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFD5,12'hFD5,12'hFD4,12'hFD4,12'hFC4,12'hFC4,12'hEC4,12'hED4,12'hEC4,12'hEC4,12'hFC4,12'hFD4,12'hEC4,12'hEC5,12'hEC4,12'hED4,12'hED4,12'hFC4,12'hED4,12'hED4,12'hFD4,12'hFD4,12'hFD5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFD4,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hEC2,12'hEB1,12'hDB3,12'hFFD,12'hFFC,12'hACB,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hBDE,12'hCC9,12'hFFE,12'hFD7,12'hED7,12'hFEA,12'hFFC,12'hFFB,12'hFE9,12'hFD6,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFD5,12'hFD5,12'hFD5,12'hFD4,12'hED4,12'hEC4,12'hFC4,12'hFC4,12'hFC4,12'hFD4,12'hFD4,12'hFD4,12'hFD5,12'hFD5,12'hFE5,12'hFD5,12'hFE5,12'hFE5,12'hFE4,12'hFE4,12'hFE4,12'hFD4,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hEB1,12'hEB2,12'hFEA,12'hFFE,12'hAB9,12'hADF,12'hAEF,
        12'hAEF,12'hAEF,12'hBDD,12'hFFD,12'hFFD,12'hED6,12'hFFC,12'hFEA,12'hFE7,12'hEE6,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFD5,12'hFD5,12'hFD5,12'hFE5,12'hFD5,12'hFE5,12'hFD5,12'hFD5,12'hFE5,12'hFE5,12'hFE5,12'hFE4,12'hFE4,12'hFD4,12'hFD4,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hEC2,12'hEB1,12'hEC6,12'hFFF,12'hAA7,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hBDC,12'hFFD,12'hFFC,12'hED6,12'hFFE,12'hFE8,12'hFD5,12'hFD5,12'hFE5,12'hFD5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFD5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFD5,12'hDB3,12'hFD4,12'hFE5,12'hFE4,12'hFD4,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hEB1,12'hDB5,12'hFFE,12'hAA7,12'h9EF,12'hADF,
        12'hAEF,12'hAEF,12'hBCB,12'hFFE,12'hFFC,12'hED7,12'hFE9,12'hFE6,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hDB3,12'hDC4,12'hDC4,12'hFD4,12'hFD4,12'hFD5,12'hFE5,12'hFD4,12'hEC4,12'hEC4,12'hFD4,12'hFE5,12'hFE5,12'hFE5,12'hFD5,12'hEC4,12'hFF9,12'hDB3,12'hFD4,12'hFD4,12'hFD4,12'hFD3,12'hFD3,12'hED3,12'hFD2,12'hFD3,12'hFD3,12'hFD3,12'hEB2,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hEB2,12'hDB4,12'hFFE,12'hCB9,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAB9,12'hFFE,12'hFEB,12'hFE7,12'hED6,12'hFE5,12'hFE4,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFD5,12'hED6,12'hFFB,12'hFEA,12'hEC7,12'hDB4,12'hFD5,12'hFE5,12'hDB3,12'hEE8,12'hED8,12'hCB3,12'hFD5,12'hFE5,12'hFE4,12'hFD4,12'hDB4,12'hFFC,12'hDC6,12'hFD4,12'hFD3,12'hFD3,12'hFD3,12'hDB3,12'hDC5,12'hEC3,12'hFD3,12'hFD3,12'hDB5,12'hFD6,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hEB2,12'hDB3,12'hFFE,12'hDDA,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAB9,12'hFFE,12'hFEB,12'hEC4,12'hFD4,12'hFE5,12'hFE4,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hED8,12'hFFF,12'hFFE,12'hFFD,12'hFEB,12'hDB4,12'hFE5,12'hDB4,12'hFFC,12'hFFD,12'hCB4,12'hFD4,12'hFE4,12'hFD4,12'hFD4,12'hEC7,12'hFFE,12'hFFB,12'hEC4,12'hFD3,12'hFD3,12'hFD3,12'hDB4,12'hFFC,12'hEC6,12'hFD3,12'hDB3,12'hFFC,12'hFEA,12'hFD4,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hEB2,12'hEB3,12'hFFE,12'hEDB,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hABA,12'hFFE,12'hFEA,12'hEC4,12'hED4,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFD5,12'hED8,12'hFFE,12'hFFD,12'hFFD,12'hFFE,12'hEC6,12'hFD5,12'hDB4,12'hFFD,12'hFFE,12'hCB4,12'hFD3,12'hFD3,12'hFD3,12'hEC3,12'hFFB,12'hFFE,12'hFFD,12'hDB4,12'hFD3,12'hFD3,12'hFD3,12'hDC6,12'hFFE,12'hFFC,12'hCB4,12'hFE9,12'hFFE,12'hFFB,12'hEC3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hEB2,12'hEB2,12'hFFE,12'hEDB,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hBBA,12'hFFF,12'hFFA,12'hFC4,12'hED4,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hED8,12'hFFE,12'hFEB,12'hFEB,12'hFFE,12'hFE9,12'hFD5,12'hDB3,12'hFFD,12'hFFE,12'hCB4,12'hFD3,12'hFD3,12'hFD3,12'hDB3,12'hFFC,12'hFFE,12'hFFE,12'hED8,12'hFD3,12'hFD3,12'hFD3,12'hFE9,12'hFFE,12'hFFE,12'hDD8,12'hFFC,12'hFFE,12'hED7,12'hEC3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hEB1,12'hEB2,12'hFFE,12'hEDB,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAB9,12'hFFF,12'hFFA,12'hFC4,12'hED4,12'hFD5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hED8,12'hFFE,12'hFFB,12'hFEA,12'hFFE,12'hFEA,12'hFD4,12'hDB3,12'hFFD,12'hFFE,12'hCB3,12'hFD3,12'hFD3,12'hFD3,12'hEC7,12'hFFE,12'hFEB,12'hFFE,12'hFFC,12'hDC3,12'hFD3,12'hFD3,12'hCB3,12'hFFB,12'hFFE,12'hFFD,12'hFFD,12'hFEA,12'hDC3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFC2,12'hEB2,12'hEB2,12'hFFE,12'hEDB,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'h9B9,12'hFFE,12'hFFB,12'hFC4,12'hFC4,12'hFD4,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hED8,12'hFFE,12'hFFB,12'hFFB,12'hFFE,12'hFD8,12'hFD3,12'hDB3,12'hFFD,12'hFFE,12'hCB3,12'hFD3,12'hFD3,12'hEC3,12'hFFB,12'hFFE,12'hCB5,12'hFFD,12'hFFD,12'hDB5,12'hFD3,12'hFD3,12'hFD3,12'hCB4,12'hFFD,12'hFFF,12'hFFC,12'hCB4,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hEB1,12'hEB2,12'hDB3,12'hFFE,12'hDCA,12'hAEF,12'hAEF,
        12'h9EF,12'hAEF,12'hBDC,12'hFFE,12'hFFC,12'hFD4,12'hEC4,12'hFC4,12'hFD4,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFD5,12'hED8,12'hFFE,12'hFFD,12'hFFD,12'hFFD,12'hDA3,12'hFD3,12'hDB3,12'hFFD,12'hFFE,12'hCB3,12'hFD3,12'hFD3,12'hCB4,12'hFFD,12'hFFD,12'hCA4,12'hFFC,12'hFFE,12'hFEA,12'hED3,12'hFD3,12'hFD3,12'hEC4,12'hFFB,12'hFFE,12'hFFB,12'hEC3,12'hFD3,12'hFD4,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hEB1,12'hEB1,12'hDB4,12'hFFE,12'hCB8,12'hAEF,12'hAEF,
        12'h9EF,12'hAEF,12'hBED,12'hFED,12'hFFD,12'hFD4,12'hEC5,12'hFC4,12'hFC4,12'hFD5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hFE5,12'hED8,12'hFFE,12'hFFE,12'hFFD,12'hEE9,12'hFC4,12'hFD3,12'hDB3,12'hFFD,12'hFFE,12'hCB4,12'hFD3,12'hFD3,12'hED7,12'hFFE,12'hFFE,12'hFEA,12'hFFD,12'hFFE,12'hFFD,12'hCB3,12'hFD2,12'hFD3,12'hFD3,12'hED9,12'hFFE,12'hFEB,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hEB1,12'hEB1,12'hEB1,12'hEB5,12'hFFF,12'hA97,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hBDE,12'hCC9,12'hFFE,12'hFD6,12'hFC4,12'hFC4,12'hFC4,12'hEC4,12'hFD5,12'hFE5,12'hFE5,12'hFD5,12'hFE5,12'hFE5,12'hFE5,12'hED8,12'hFFE,12'hFFD,12'hED7,12'hDB3,12'hFD3,12'hFD3,12'hDB3,12'hFFD,12'hFFE,12'hDB3,12'hFD3,12'hEC3,12'hFFB,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hEC7,12'hFD3,12'hFD3,12'hFD4,12'hEC7,12'hFFE,12'hFE9,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD4,12'hFD3,12'hEB2,12'hEB2,12'hEB1,12'hEB2,12'hEC7,12'hFFE,12'hAA9,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hBEF,12'hAA7,12'hFFF,12'hFE7,12'hFC4,12'hFC4,12'hFC4,12'hEC4,12'hEC4,12'hFD4,12'hFD5,12'hFE5,12'hFE5,12'hFE5,12'hFD5,12'hED8,12'hFFE,12'hFEB,12'hEC4,12'hFD3,12'hFD3,12'hFD3,12'hDB3,12'hFFD,12'hFFE,12'hCB4,12'hFD3,12'hDB3,12'hFFD,12'hFFE,12'hFFC,12'hFFB,12'hFEA,12'hFFD,12'hFFE,12'hFF9,12'hEC3,12'hFD3,12'hFD3,12'hEC6,12'hFFF,12'hFE9,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hFC2,12'hEB2,12'hDC5,12'hFE9,12'hDB3,12'hEB2,12'hFEB,12'hFFE,12'hABA,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'h9A8,12'hFFF,12'hFFA,12'hEC5,12'hFC4,12'hFC4,12'hEC4,12'hFC4,12'hFC4,12'hFC4,12'hED4,12'hFD5,12'hFE5,12'hFD5,12'hED8,12'hFFE,12'hFE9,12'hFD3,12'hFD3,12'hFD3,12'hFD3,12'hDB3,12'hFFE,12'hFFE,12'hED9,12'hED6,12'hDB4,12'hFFB,12'hFFC,12'hCB4,12'hDB3,12'hDB3,12'hEE9,12'hFFC,12'hDB5,12'hFD3,12'hFD3,12'hFD3,12'hED6,12'hFFE,12'hFE9,12'hFD3,12'hFD3,12'hFD3,12'hEC2,12'hEB2,12'hEB1,12'hDB3,12'hFFB,12'hFFD,12'hED8,12'hDB3,12'hFFD,12'hFFC,12'hBCB,12'hAEF,12'hAEF,
        12'hAEF,12'hAEE,12'hAEF,12'hACB,12'hFFC,12'hFFE,12'hFD5,12'hFC4,12'hFC4,12'hEC4,12'hFC4,12'hFC4,12'hFC4,12'hFD4,12'hFC4,12'hFC4,12'hEB3,12'hDB3,12'hED8,12'hFE7,12'hEC2,12'hFC3,12'hFD3,12'hFD3,12'hDB3,12'hFFD,12'hFFE,12'hFFE,12'hFFD,12'hDB4,12'hDB4,12'hFE7,12'hED4,12'hFD3,12'hFD3,12'hDB3,12'hDB5,12'hFD4,12'hFD3,12'hFC2,12'hFC3,12'hEC5,12'hFFB,12'hFD7,12'hEB2,12'hEB2,12'hEB1,12'hEB1,12'hEB2,12'hEB1,12'hEC6,12'hFFD,12'hFFE,12'hFFA,12'hDB5,12'hFFE,12'hDC9,12'hBDE,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hBDE,12'hCC8,12'hFFF,12'hEE8,12'hEC4,12'hFC4,12'hED3,12'hFC4,12'hFC4,12'hFC4,12'hFC4,12'hFC4,12'hEB3,12'hEB2,12'hEB1,12'hEB2,12'hDB2,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hDB2,12'hFFA,12'hFFC,12'hFFC,12'hFFC,12'hCA3,12'hEB2,12'hDB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB1,12'hEB1,12'hEB2,12'hDA2,12'hDA3,12'hDB2,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hFFB,12'hFFE,12'hFFE,12'hFFB,12'hEEA,12'hFFF,12'hA96,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'h9A6,12'hFFE,12'hFFC,12'hED5,12'hFC4,12'hFC4,12'hFC4,12'hFC4,12'hEC4,12'hFC4,12'hEC3,12'hEB2,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB2,12'hEB1,12'hEB2,12'hDB3,12'hDA4,12'hDB4,12'hDB5,12'hDB3,12'hEB1,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hEB1,12'hEB2,12'hEB1,12'hEB1,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB3,12'hFFD,12'hFFE,12'hFFE,12'hEDA,12'hFFE,12'hFFC,12'hBCB,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBDD,12'hEEA,12'hFFE,12'hFE9,12'hFD4,12'hFC4,12'hFC4,12'hFC4,12'hFC4,12'hFC4,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB1,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB1,12'hEB2,12'hEB2,12'hEB1,12'hEB1,12'hEB1,12'hEB2,12'hDB5,12'hFFE,12'hFFE,12'hFFD,12'hEDB,12'hFFF,12'hBB6,12'hADF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hADF,12'h9A6,12'hFFF,12'hFFE,12'hFE7,12'hEC4,12'hFC4,12'hFC4,12'hFD4,12'hEB2,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB2,12'hEB1,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB1,12'hEB1,12'hEB2,12'hEB2,12'hEB1,12'hEB2,12'hDB3,12'hFE8,12'hED8,12'hFFB,12'hFFC,12'hDDA,12'hFFD,12'hFFD,12'hAB9,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'h9EF,12'hCDE,12'hCB8,12'hFFF,12'hFFC,12'hFD7,12'hFD4,12'hFC4,12'hEC3,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB1,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB2,12'hEB2,12'hEB1,12'hEB2,12'hEB1,12'hEB1,12'hEB2,12'hEB1,12'hEB2,12'hDB5,12'hFFD,12'hFFA,12'hDB4,12'hCB5,12'hFFD,12'hFFF,12'hAA6,12'hBDE,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hADF,12'hABB,12'hEDB,12'hFFE,12'hFFC,12'hFD8,12'hFC4,12'hDB2,12'hEB2,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB2,12'hEB1,12'hEB1,12'hEB1,12'hEB2,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB1,12'hEB2,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hEB3,12'hFE6,12'hFE8,12'hDB5,12'hEC4,12'hFFB,12'hFFF,12'hDD9,12'hBCB,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hADE,12'hAA7,12'hFEB,12'hFFF,12'hFFD,12'hFE9,12'hFD5,12'hEC3,12'hEB3,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB2,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB1,12'hEB2,12'hEB1,12'hEB1,12'hEB2,12'hEB1,12'hEB1,12'hEB2,12'hEB4,12'hEC5,12'hEE8,12'hFFD,12'hFFF,12'hEEB,12'hAB9,12'hADF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBDE,12'h9A8,12'hEDA,12'hFFE,12'hFFE,12'hFFE,12'hFFB,12'hFE9,12'hFE8,12'hFE7,12'hED6,12'hED6,12'hFD5,12'hEC5,12'hEC4,12'hEC3,12'hEC3,12'hEC3,12'hEC2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB3,12'hEC3,12'hEC3,12'hEC3,12'hEC4,12'hEC4,12'hEC4,12'hED5,12'hED5,12'hED6,12'hFD7,12'hFD7,12'hFE8,12'hFEA,12'hFFD,12'hFFE,12'hFFF,12'hEEB,12'hAA9,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAB9,12'hBB8,12'hFEC,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFD,12'hFFD,12'hFFC,12'hFFC,12'hFFB,12'hFFA,12'hFEA,12'hFE9,12'hFE8,12'hFE8,12'hFE8,12'hFE8,12'hFE8,12'hFE8,12'hFE8,12'hFE8,12'hFE9,12'hFEA,12'hFFA,12'hFFB,12'hFFB,12'hFFB,12'hFFC,12'hFFC,12'hFFD,12'hFFD,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFF,12'hFFD,12'hCB8,12'hAB9,12'hBDF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hADC,12'hAA8,12'hAA6,12'hCC9,12'hFEC,12'hFFD,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hEDB,12'hBB8,12'h9A7,12'hBCB,12'hADF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hADF,12'hBEF,12'hBDE,12'hBDD,12'hABA,12'h9A9,12'hAA7,12'hA97,12'hAA7,12'hBA8,12'hBB8,12'hCC9,12'hDDA,12'hDDA,12'hEDA,12'hEEB,12'hEEC,12'hFEC,12'hFFC,12'hFFD,12'hFFC,12'hFED,12'hFEC,12'hFEC,12'hEEC,12'hEEB,12'hEDA,12'hDDA,12'hDDA,12'hDC9,12'hCB8,12'hBA7,12'hBA7,12'hAA7,12'h9A7,12'h9B8,12'h9B9,12'hACB,12'hBDD,12'hBDE,12'hADF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEE,12'hADE,12'hBDE,12'hBDD,12'hABB,12'hBCA,12'hBB9,12'hAA8,12'hAB8,12'hAA8,12'hAA8,12'hAA8,12'hAA8,12'hAB8,12'hAA8,12'hAA8,12'hBCB,12'hBCC,12'hACB,12'hBEE,12'hBED,12'hBDD,12'hAEE,12'hAEF,12'hAEF,12'hAEF,12'hADF,12'hADF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hADF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hADF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF

    };


    always @(*) begin
        if(h_cnt >= 290 && h_cnt <= 349 && v_cnt >= 335 && v_cnt <= 374) begin
            if(play[(v_cnt - 335) * 60 + (h_cnt - 290)] != 12'hAEF) begin
                background = 0;
                vga = play[(v_cnt - 335) * 60 + (h_cnt - 290)];
            end
            else begin
                background = 1;
                vga = 12'h000;
            end
        end
        else begin
            background = 1;
            vga = 12'h000;
        end
    end
endmodule

module reverse (
    input [9:0] h_cnt,
    input [9:0] v_cnt,
    output reg background, //1 for print background 0 for print fish
    output reg [11:0] vga
);
    parameter [11:0] reverse [0:719] = {//24*30
  
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBDD,12'hAB9,12'hAB8,12'hAB8,12'hBB8,12'hBCD,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBEE,12'hABA,12'hBA6,12'hDCA,12'hFFC,12'hFFE,12'hFFE,12'hFFE,12'hEEA,12'hAA6,12'hAA8,12'hBDE,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBDE,12'hA97,12'hFEB,12'hFFE,12'hFFE,12'hFFE,12'hFFD,12'hFFE,12'hFFE,12'hFFF,12'hFFF,12'hFFD,12'hBA7,12'hBCB,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBDD,12'hBA7,12'hFFD,12'hFFE,12'hFFB,12'hDC6,12'hEB4,12'hDB3,12'hDB3,12'hDB3,12'hDC6,12'hFEA,12'hFFE,12'hFFF,12'hDD9,12'hBBA,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBA6,12'hFFE,12'hFFE,12'hDC7,12'hEB3,12'hEB1,12'hEB2,12'hEB2,12'hEB1,12'hEB2,12'hEB1,12'hEB3,12'hDB4,12'hFFC,12'hFFF,12'hDDA,12'hBDC,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAA6,12'hFFF,12'hFFE,12'hDC8,12'hFE9,12'hEC4,12'hEC2,12'hFC3,12'hEC3,12'hFC3,12'hFC3,12'hFC3,12'hFC2,12'hEB2,12'hDB2,12'hFEC,12'hFFF,12'hCB8,12'hBEE,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hBCB,12'hFFB,12'hFFE,12'hDD7,12'hFFD,12'hFFE,12'hFFA,12'hEC3,12'hFC3,12'hFC2,12'hFC3,12'hEC2,12'hFD2,12'hFC2,12'hFC3,12'hEB2,12'hDB3,12'hFFC,12'hFFE,12'hB96,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hBA7,12'hFFF,12'hFE9,12'hDC7,12'hFFD,12'hFFB,12'hFD5,12'hFC2,12'hEC3,12'hDB3,12'hEB3,12'hEC3,12'hFD3,12'hFC2,12'hFC2,12'hFC3,12'hEB2,12'hEB5,12'hFFE,12'hFEB,12'hBCC,12'hAEF,
        12'hAEF,12'hBCA,12'hFFD,12'hFFD,12'hDC5,12'hFEA,12'hED5,12'hFC4,12'hEC2,12'hDB5,12'hFE9,12'hFFB,12'hFFB,12'hED8,12'hCB4,12'hEC3,12'hFC2,12'hFC2,12'hFC3,12'hEB2,12'hFEA,12'hFFE,12'hA96,12'hAEF,
        12'hAEF,12'h995,12'hFFF,12'hFE8,12'hEC4,12'hED5,12'hFC2,12'hDB3,12'hED9,12'hFFD,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFC,12'hDC7,12'hEC3,12'hFC3,12'hEC2,12'hEC2,12'hDB4,12'hFFF,12'hDD9,12'hBDE,
        12'hBEE,12'hCC8,12'hFFF,12'hEC5,12'hEC3,12'hFC3,12'hEC3,12'hED9,12'hFFE,12'hFFE,12'hFFF,12'hFFE,12'hFFD,12'hFFE,12'hFFE,12'hFFD,12'hDB4,12'hFC3,12'hFC3,12'hFC3,12'hDB2,12'hFFC,12'hFFD,12'hBCA,
        12'hBDC,12'hFFC,12'hFFD,12'hEC3,12'hFC2,12'hFC3,12'hDB4,12'hFFD,12'hFFE,12'hFFE,12'hFFB,12'hFD9,12'hED9,12'hFFD,12'hFFE,12'hFFE,12'hFFC,12'hDB3,12'hFC2,12'hEC3,12'hEB2,12'hED8,12'hFFE,12'hAA8,
        12'hAB9,12'hFFE,12'hFEA,12'hEB1,12'hFC2,12'hFC3,12'hFEA,12'hFFE,12'hFFE,12'hFEA,12'hDB3,12'hEC2,12'hEC3,12'hDB4,12'hFFC,12'hFFE,12'hFFE,12'hDC6,12'hFC2,12'hED2,12'hFC2,12'hDB4,12'hFFF,12'hA96,
        12'hABA,12'hFFF,12'hFE8,12'hEB2,12'hED2,12'hDB3,12'hFFD,12'hFFE,12'hFFD,12'hDB3,12'hFC3,12'hFC2,12'hEC3,12'hDB4,12'hDC8,12'hFFE,12'hFFE,12'hFEB,12'hDB3,12'hEC3,12'hFC3,12'hDB4,12'hFFF,12'hBA7,
        12'hABA,12'hFFE,12'hFE7,12'hEB2,12'hFC2,12'hDB3,12'hFFE,12'hFFE,12'hFEA,12'hEB2,12'hEB2,12'hEB2,12'hEC5,12'hFFC,12'hFFD,12'hFFE,12'hFFE,12'hFFD,12'hFFC,12'hEC5,12'hFC3,12'hDB3,12'hFFE,12'hDC8,
        12'hABA,12'hFFF,12'hFD7,12'hEB2,12'hFC2,12'hDB4,12'hFFE,12'hFFE,12'hED7,12'hEB1,12'hEB1,12'hEB2,12'hFE9,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFEA,12'hFC3,12'hDB3,12'hFFE,12'hDC9,
        12'hABA,12'hFFF,12'hFE8,12'hEB2,12'hFC2,12'hDB3,12'hFFE,12'hFFE,12'hED8,12'hEB1,12'hEB2,12'hEB2,12'hDC6,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFD,12'hEC7,12'hFC3,12'hDB3,12'hFFE,12'hCB8,
        12'hAB9,12'hFFE,12'hFE9,12'hEB1,12'hFC2,12'hDA2,12'hFFD,12'hFFE,12'hFFB,12'hDB2,12'hEB2,12'hEB2,12'hDA3,12'hFFC,12'hFFE,12'hFFE,12'hFFE,12'hFFF,12'hFFD,12'hDA3,12'hFC2,12'hDB4,12'hFFF,12'hA96,
        12'hADC,12'hFFD,12'hFFB,12'hEB2,12'hEB2,12'hEB2,12'hFFC,12'hFFE,12'hFFE,12'hDC6,12'hEB2,12'hEB2,12'hEB2,12'hDC6,12'hFFD,12'hFFE,12'hFFE,12'hFFD,12'hEC7,12'hEB2,12'hEB1,12'hEC7,12'hFFF,12'hA97,
        12'hBDE,12'hED9,12'hFFD,12'hEC4,12'hEB2,12'hEB2,12'hED7,12'hFFE,12'hFFE,12'hFFD,12'hED7,12'hDB3,12'hEB1,12'hEB2,12'hED8,12'hFFD,12'hFFD,12'hFD8,12'hDB4,12'hED7,12'hEB3,12'hFEB,12'hFFE,12'hAB9,
        12'hAEF,12'hBA6,12'hFFF,12'hED7,12'hEB1,12'hEB1,12'hDB3,12'hFFC,12'hFFE,12'hFFE,12'hFFD,12'hFFB,12'hDB3,12'hEB1,12'hEB2,12'hDB4,12'hDB4,12'hDB3,12'hFFC,12'hFFD,12'hDB5,12'hFFE,12'hEEB,12'hBED,
        12'hAEF,12'h9BA,12'hFFE,12'hFFC,12'hEC3,12'hEB2,12'hEB2,12'hDB4,12'hFFD,12'hFFE,12'hFFF,12'hFFD,12'hDB3,12'hEB1,12'hEB2,12'hEB2,12'hEB1,12'hEB4,12'hFFD,12'hFFD,12'hED8,12'hFFF,12'hB97,12'hAEF,
        12'hAEF,12'hBDD,12'hCC9,12'hFFF,12'hED7,12'hEB2,12'hEB2,12'hEB2,12'hDB4,12'hFFB,12'hFFC,12'hFFB,12'hDB2,12'hEB1,12'hEB2,12'hEB1,12'hEB3,12'hDC6,12'hFFD,12'hFEA,12'hFFE,12'hFFD,12'hBBA,12'hAEF,
        12'hAEF,12'hAEF,12'hAB8,12'hFFD,12'hFFD,12'hFD5,12'hEB1,12'hEB2,12'hEB1,12'hDB3,12'hDB4,12'hDB3,12'hEB2,12'hEB1,12'hEB1,12'hEB2,12'hFD7,12'hFE9,12'hDB5,12'hEEA,12'hFFF,12'hAA7,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hBA7,12'hFFF,12'hFFC,12'hED4,12'hEB1,12'hEB1,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hDB3,12'hEB3,12'hFD8,12'hFFF,12'hEDB,12'hBCB,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hBDD,12'hDD9,12'hFFF,12'hFFC,12'hED6,12'hEC2,12'hEB2,12'hEB1,12'hEB2,12'hEB1,12'hEB2,12'hEB1,12'hEB2,12'hEC3,12'hFE9,12'hFFF,12'hFFC,12'hAA8,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBDC,12'hEC9,12'hFFE,12'hFFD,12'hFE9,12'hED5,12'hEC3,12'hEB2,12'hEB2,12'hEB3,12'hEC4,12'hED8,12'hFFC,12'hFFF,12'hFFD,12'hA97,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBCA,12'hBB8,12'hFFD,12'hFFE,12'hFFD,12'hFFC,12'hFEA,12'hFFA,12'hFFB,12'hFFD,12'hFFE,12'hFFF,12'hEDA,12'hAA8,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBDD,12'h997,12'hCC9,12'hFFE,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFD,12'hEDA,12'hA95,12'hACB,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBDD,12'hAB9,12'hAA6,12'hAA7,12'hBB7,12'hAA6,12'hAA8,12'hBDC,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF

    };


    always @(*) begin
        if(h_cnt >= 308 && h_cnt <= 331 && v_cnt >= 340 && v_cnt <= 369) begin
            if(reverse[(v_cnt - 340) * 24 + (h_cnt - 308)] != 12'hAEF) begin
                background = 0;
                vga = reverse[(v_cnt - 340) * 24 + (h_cnt - 308)];
            end
            else begin
                background = 1;
                vga = 12'h000;
            end
        end
        else begin
            background = 1;
            vga = 12'h000;
        end
    end
endmodule

module pause (
    input [9:0] h_cnt,
    input [9:0] v_cnt,
    input pause_in,
    output reg background, //1 for print background 0 for print fish
    output reg [11:0] vga
);
    parameter [11:0] pause1 [0:719] = {//24*30
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hADC,12'hBCC,12'hBDC,12'hADC,12'hBDD,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hACB,12'hAA8,12'hCB8,12'hEDB,12'hFFD,12'hFFD,12'hFEC,12'hDC9,12'hAA7,12'hAB9,12'hBEE,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'h9EE,12'hAEF,12'hAEF,12'h9A7,12'hDD9,12'hFFF,12'hFFF,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFF,12'hFFF,12'hFFC,12'hBA7,12'hBDC,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hA95,12'hFFD,12'hFFF,12'hFFD,12'hED9,12'hDB5,12'hDB4,12'hDB3,12'hDB4,12'hEC6,12'hFEA,12'hFFF,12'hFFE,12'hDD9,12'hBBB,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBA6,12'hFFE,12'hFFE,12'hED9,12'hDB3,12'hEB2,12'hEB1,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hEB3,12'hDC5,12'hFFC,12'hFFF,12'hEEB,12'hBCA,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'h9A7,12'hFFE,12'hFFE,12'hDC9,12'hFD8,12'hDB4,12'hFC2,12'hFC3,12'hFC2,12'hFC2,12'hFC3,12'hFC2,12'hEC2,12'hEB1,12'hDB3,12'hFEB,12'hFFF,12'hDCA,12'hADD,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hACB,12'hFFD,12'hFFE,12'hDC8,12'hFFC,12'hFFD,12'hFE9,12'hED3,12'hFC3,12'hFC2,12'hFC2,12'hEC3,12'hFC2,12'hFC2,12'hFC2,12'hEB2,12'hDB3,12'hFFB,12'hFFE,12'hAA6,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hBB7,12'hFFF,12'hFE9,12'hEC7,12'hFFD,12'hFFD,12'hED7,12'hED3,12'hEC3,12'hFC3,12'hFC2,12'hFC2,12'hFC3,12'hFC3,12'hFC2,12'hFC2,12'hEB2,12'hDB4,12'hFFE,12'hFFD,12'hABA,12'hAEF,
        12'hAEF,12'hABA,12'hFFD,12'hFFD,12'hDC5,12'hFEA,12'hFE7,12'hEC4,12'hEC2,12'hDB5,12'hFFA,12'hFEA,12'hCB4,12'hEC3,12'hEC2,12'hFC2,12'hFC2,12'hFC2,12'hFC3,12'hEB1,12'hED8,12'hFFE,12'hBA7,12'hAEF,
        12'hAEF,12'hB97,12'hFFF,12'hFE8,12'hEC5,12'hEE7,12'hED3,12'hFC2,12'hDB3,12'hFFC,12'hFFE,12'hFFE,12'hFFE,12'hFD8,12'hDB3,12'hFC3,12'hFC2,12'hFC2,12'hEC2,12'hFC3,12'hDB4,12'hFFD,12'hFFB,12'hBDC,
        12'hBDD,12'hDDA,12'hFFE,12'hEC4,12'hFC4,12'hEC2,12'hEC3,12'hFC2,12'hDB5,12'hFFD,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFEA,12'hDB3,12'hFC2,12'hFC3,12'hFC3,12'hFC2,12'hEB2,12'hFD9,12'hFFF,12'hAA7,
        12'hBDC,12'hFFD,12'hFFC,12'hEB2,12'hFC3,12'hFC2,12'hFC3,12'hFC3,12'hED7,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFE9,12'hEC3,12'hFC2,12'hEC3,12'hFC2,12'hEC2,12'hDB4,12'hFFF,12'hAA6,
        12'h9A8,12'hFFE,12'hFE9,12'hEB2,12'hFC2,12'hFC2,12'hFC3,12'hFC3,12'hFE9,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFD,12'hDC6,12'hFC3,12'hFC2,12'hFC2,12'hFC2,12'hDB3,12'hFFE,12'hDCA,
        12'hAA7,12'hFFE,12'hED7,12'hEB2,12'hFC2,12'hFC2,12'hFC2,12'hFC3,12'hFE9,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFC,12'hDB3,12'hFC2,12'hFC3,12'hFC3,12'hEB3,12'hFFD,12'hEEC,
        12'hAA7,12'hFFF,12'hED6,12'hEC2,12'hFC2,12'hFC3,12'hFC3,12'hFC3,12'hFEA,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFD,12'hDB4,12'hFC3,12'hEC3,12'hFC3,12'hEB2,12'hFFD,12'hFFD,
        12'hAA7,12'hFFF,12'hFD5,12'hEC2,12'hFC2,12'hED3,12'hFC3,12'hFC2,12'hFEA,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hED7,12'hFC3,12'hFC3,12'hFC3,12'hEB2,12'hFFC,12'hFFD,
        12'hAA6,12'hFFF,12'hFD6,12'hEC2,12'hFC2,12'hFC3,12'hEC2,12'hEB2,12'hFEA,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hDC5,12'hFC2,12'hFC3,12'hFC3,12'hEB2,12'hFFD,12'hFFD,
        12'h9A8,12'hFFF,12'hFE8,12'hDB2,12'hFC3,12'hEB1,12'hEB2,12'hEB2,12'hFE9,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFC,12'hDB3,12'hEB1,12'hEC1,12'hEC2,12'hDB3,12'hFFD,12'hDEB,
        12'hAB9,12'hFFE,12'hFEA,12'hDB2,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hFD9,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hED8,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hDB3,12'hFFE,12'hBB9,
        12'hBDC,12'hFFC,12'hFFD,12'hEC3,12'hEB2,12'hEB2,12'hEB2,12'hFB2,12'hFD8,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFC,12'hDB2,12'hEB2,12'hEB3,12'hFD6,12'hEB2,12'hEC6,12'hFFF,12'h997,
        12'hBEE,12'hCC8,12'hFFE,12'hED6,12'hEB2,12'hEB1,12'hEB2,12'hEB1,12'hDC6,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFE,12'hFFC,12'hCB4,12'hEB1,12'hEB2,12'hFE8,12'hFFD,12'hDC5,12'hFEB,12'hFFE,12'hAB9,
        12'hAEF,12'hAA7,12'hFFE,12'hFFA,12'hEB3,12'hEB1,12'hEB2,12'hEB2,12'hDB2,12'hFFD,12'hFFE,12'hFFE,12'hFFD,12'hFFC,12'hDB4,12'hEB2,12'hEB1,12'hDB3,12'hFFD,12'hFFE,12'hDC8,12'hFFE,12'hDD9,12'hBDD,
        12'hAEF,12'hBDD,12'hFEB,12'hFFE,12'hED6,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hFD8,12'hFFD,12'hFFD,12'hFE9,12'hDB3,12'hEB1,12'hEB1,12'hEB2,12'hDB4,12'hFFD,12'hFFC,12'hFFC,12'hFFF,12'h998,12'hAEF,
        12'hAEF,12'hAEF,12'hAA7,12'hFFF,12'hFFC,12'hEC4,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hDB4,12'hDB3,12'hDB2,12'hEB1,12'hEB2,12'hEB2,12'hEC5,12'hFF9,12'hDC5,12'hDC8,12'hFFE,12'hDDA,12'hBDC,12'hAEF,
        12'hAEF,12'hAEF,12'hBDD,12'hCC9,12'hFFF,12'hFFB,12'hEC4,12'hEB2,12'hEB1,12'hEB1,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEC4,12'hDB4,12'hDC5,12'hFFE,12'hFFE,12'hAA7,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hBCA,12'hEEB,12'hFFF,12'hFFB,12'hED5,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEC7,12'hFFD,12'hFFE,12'hAA7,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAB9,12'hFEB,12'hFFE,12'hFFD,12'hFE8,12'hED4,12'hEC2,12'hEB2,12'hEB1,12'hEB2,12'hEC3,12'hFD6,12'hFFA,12'hFFE,12'hFFE,12'hA96,12'hBDD,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBB9,12'hDCA,12'hFFE,12'hFFF,12'hFFE,12'hFFB,12'hFEA,12'hFEA,12'hFFB,12'hFFC,12'hFFE,12'hFFF,12'hFFC,12'hA97,12'hADD,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBDC,12'hA96,12'hEDA,12'hFFD,12'hFFF,12'hFFF,12'hFFF,12'hFFE,12'hFFF,12'hFFD,12'hBB6,12'hAB9,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBDC,12'hABA,12'hAA7,12'hAA7,12'hBB8,12'hBA7,12'hAA7,12'hACB,12'hBDE,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF
        
    };

    parameter [11:0] pause2 [0:719] = {//24*30
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBDD,12'hACC,12'hACB,12'hBCD,12'hBDE,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBDC,12'hAB7,12'hBA7,12'hDCA,12'hEEC,12'hEEB,12'hDDA,12'hBB8,12'hAA7,12'hACA,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBDE,12'hAB8,12'hCC8,12'hFFE,12'hFFF,12'hFFF,12'hFFF,12'hFFE,12'hFFE,12'hFFF,12'hFFF,12'hEEC,12'hA96,12'hBDC,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hBDD,12'h9A7,12'hFFD,12'hFFF,12'hFFD,12'hFEA,12'hEC6,12'hEB4,12'hDB4,12'hDB5,12'hED7,12'hFFB,12'hFFE,12'hFFE,12'hCB9,12'hBDC,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'h997,12'hFFE,12'hFFE,12'hFEA,12'hDB4,12'hEB2,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hDB2,12'hEC6,12'hFFD,12'hFFE,12'hEDA,12'hBCB,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'h9A8,12'hFFD,12'hFFF,12'hDD9,12'hDC6,12'hDB3,12'hEC2,12'hFC2,12'hFC2,12'hFC2,12'hFC2,12'hFC2,12'hEC2,12'hEB2,12'hDB3,12'hFFC,12'hFFE,12'hCB9,12'hBDD,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hBDC,12'hFEC,12'hFFE,12'hED9,12'hFFC,12'hFFE,12'hFF9,12'hFC3,12'hFC2,12'hED2,12'hFC2,12'hFC2,12'hFC2,12'hEC2,12'hFC3,12'hEB2,12'hDB3,12'hFFD,12'hFFE,12'h9A7,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hBA7,12'hFFE,12'hFEA,12'hDD6,12'hFFD,12'hFFD,12'hFE6,12'hEC3,12'hFC2,12'hFC3,12'hFC2,12'hFC3,12'hFC3,12'hFC3,12'hFC2,12'hFC3,12'hEB2,12'hDB4,12'hFFD,12'hFFD,12'hBCA,12'hAEF,
        12'hAEF,12'hBBA,12'hFFC,12'hFFE,12'hEC5,12'hEE9,12'hFE8,12'hED5,12'hED3,12'hFC3,12'hFC2,12'hFC2,12'hFC2,12'hFC3,12'hFC3,12'hFC3,12'hFC2,12'hFC2,12'hFC3,12'hEB2,12'hED9,12'hFFE,12'hBA6,12'hAEF,
        12'hAEF,12'h9A7,12'hFFF,12'hFE8,12'hEC4,12'hFD7,12'hFC3,12'hFC3,12'hDB3,12'hCB3,12'hDB3,12'hFC3,12'hFC3,12'hDC2,12'hCB3,12'hCB3,12'hEC3,12'hFC3,12'hEC2,12'hFC2,12'hDB4,12'hFFD,12'hFFC,12'hBCC,
        12'hBDE,12'hDDA,12'hFFE,12'hED4,12'hFC5,12'hEC3,12'hEC2,12'hDB3,12'hFFC,12'hFFD,12'hFEA,12'hDB3,12'hEC3,12'hED8,12'hFFD,12'hFFC,12'hDC6,12'hFC2,12'hFC3,12'hFC3,12'hEB2,12'hFEA,12'hFFE,12'hAA8,
        12'hBDC,12'hFFE,12'hFFB,12'hEB3,12'hFD2,12'hFC2,12'hFC3,12'hFE9,12'hFFE,12'hFFE,12'hFFD,12'hDB5,12'hDB3,12'hFFD,12'hFFE,12'hFFE,12'hFFC,12'hDB3,12'hFC2,12'hEC3,12'hEB2,12'hDC5,12'hFFF,12'h9A6,
        12'h9A8,12'hFFE,12'hFE9,12'hEB2,12'hFC3,12'hFC2,12'hFC3,12'hFEA,12'hFFE,12'hFFE,12'hFFE,12'hDC6,12'hDB3,12'hFFE,12'hFFE,12'hFFE,12'hFFD,12'hDB3,12'hFC3,12'hFC3,12'hFC2,12'hDB3,12'hFFE,12'hCC9,
        12'hAA7,12'hFFE,12'hFE7,12'hEB2,12'hFC3,12'hFC2,12'hFC3,12'hFFA,12'hFFE,12'hFFE,12'hFFE,12'hEC7,12'hDB3,12'hFFE,12'hFFE,12'hFFE,12'hFFD,12'hDB3,12'hFC2,12'hFC2,12'hFC2,12'hEB2,12'hFFD,12'hEEC,
        12'hAA6,12'hFFF,12'hED6,12'hEC2,12'hFC3,12'hFC2,12'hFC3,12'hFFB,12'hFFE,12'hFFE,12'hFFE,12'hEC7,12'hCB3,12'hFFE,12'hFFE,12'hFFE,12'hFFD,12'hDB3,12'hFC2,12'hFC2,12'hFC2,12'hEB2,12'hFFD,12'hFFD,
        12'hBA7,12'hFFF,12'hFD5,12'hEB2,12'hFC3,12'hFC2,12'hFC3,12'hFFB,12'hFFE,12'hFFE,12'hFFE,12'hEC7,12'hCB3,12'hFFE,12'hFFE,12'hFFE,12'hFFD,12'hDB3,12'hFC3,12'hFC3,12'hFC3,12'hEB2,12'hFFC,12'hFFD,
        12'hAA6,12'hFFF,12'hFD6,12'hEC2,12'hFC2,12'hFC2,12'hEC3,12'hFFB,12'hFFE,12'hFFE,12'hFFE,12'hEC7,12'hCB3,12'hFFD,12'hFFE,12'hFFE,12'hFFD,12'hDB3,12'hFC2,12'hFC3,12'hFC3,12'hEB2,12'hFFD,12'hFFC,
        12'h9A7,12'hFFF,12'hFD8,12'hEB2,12'hFC3,12'hEC2,12'hEB2,12'hFFB,12'hFFE,12'hFFE,12'hFFE,12'hEC7,12'hCB3,12'hFFD,12'hFFE,12'hFFE,12'hFFD,12'hDB3,12'hEB1,12'hFC2,12'hFC2,12'hEB2,12'hFFE,12'hEDB,
        12'hABA,12'hFFE,12'hFEA,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hFFB,12'hFFE,12'hFFE,12'hFFE,12'hEC7,12'hCB3,12'hFFD,12'hFFE,12'hFFE,12'hFFD,12'hDB3,12'hEB2,12'hEB2,12'hEB2,12'hDB4,12'hFFF,12'hBB8,
        12'hBDC,12'hFFD,12'hFFC,12'hEC3,12'hEB2,12'hEB2,12'hEB2,12'hFFB,12'hFFE,12'hFFE,12'hFFE,12'hEC7,12'hDB3,12'hFFD,12'hFFE,12'hFFE,12'hFFD,12'hDB3,12'hEB3,12'hEC5,12'hEB2,12'hEC6,12'hFFF,12'h9A7,
        12'hBEE,12'hDC9,12'hFFE,12'hED6,12'hEB2,12'hEB2,12'hEB1,12'hFE9,12'hFFE,12'hFFE,12'hFFE,12'hDC6,12'hDB3,12'hFFC,12'hFFE,12'hFFE,12'hFFC,12'hDB3,12'hFD7,12'hFFC,12'hDB4,12'hFEB,12'hFFE,12'hAB9,
        12'hAEF,12'h996,12'hFFF,12'hFEA,12'hEB2,12'hEB1,12'hEB1,12'hDB4,12'hFFC,12'hFFE,12'hFFB,12'hDA2,12'hEB2,12'hFE9,12'hFFD,12'hFFD,12'hED7,12'hDB3,12'hFFC,12'hFFE,12'hDC7,12'hFFE,12'hEDB,12'hBDC,
        12'hAEF,12'hADC,12'hFEC,12'hFFE,12'hED6,12'hEB1,12'hEB2,12'hEB2,12'hDB4,12'hEC6,12'hDB3,12'hEB2,12'hEB1,12'hDA2,12'hEC5,12'hDC5,12'hDB3,12'hDB5,12'hFFD,12'hFFC,12'hFEC,12'hFFE,12'hA97,12'hAEF,
        12'hAEF,12'hAEF,12'h9A7,12'hFFE,12'hFFC,12'hFC4,12'hEB1,12'hEB1,12'hEB2,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEB2,12'hEC4,12'hFFA,12'hEC7,12'hDB7,12'hFFF,12'hFEA,12'hBCC,12'hAEF,
        12'hAEF,12'hAEF,12'hBDD,12'hDD9,12'hFFE,12'hFEA,12'hEC4,12'hEB1,12'hEB2,12'hEB2,12'hEB2,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB2,12'hEC5,12'hDC3,12'hDB4,12'hFFD,12'hFFD,12'hAA9,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hABA,12'hFEB,12'hFFF,12'hFEB,12'hFC5,12'hEB2,12'hEB1,12'hEB1,12'hEB2,12'hEB1,12'hEB1,12'hEB1,12'hEB1,12'hEB3,12'hEC6,12'hFFD,12'hFFE,12'hAA8,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAA8,12'hFEC,12'hFFE,12'hFFC,12'hFD7,12'hEC5,12'hEC3,12'hEB2,12'hEB2,12'hEB2,12'hEC3,12'hEC5,12'hFEA,12'hFFE,12'hFFE,12'hBB8,12'hBDE,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hABA,12'hDDA,12'hFFF,12'hFFE,12'hFFD,12'hFFA,12'hEE8,12'hFE8,12'hFE9,12'hFFC,12'hFFD,12'hFFF,12'hFFD,12'hAA6,12'hADD,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hACB,12'hA96,12'hEEC,12'hFFE,12'hFFF,12'hFFF,12'hFFF,12'hFFE,12'hFFE,12'hFFD,12'hCC8,12'hBA9,12'hBDE,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,
        12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hACA,12'h9A8,12'hAA7,12'hDC9,12'hDD9,12'hBB8,12'hAA8,12'hAA8,12'hBDD,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF,12'hAEF

        
    };


    always @(*) begin
        if(pause_in == 1'b1) begin
            if(h_cnt >= 600 && h_cnt <= 623 && v_cnt >= 10 && v_cnt <= 39) begin
                if(pause1[(v_cnt - 10) * 24 + (h_cnt - 600)] != 12'hAEF) begin
                    background = 0;
                    vga = pause1[(v_cnt - 10) * 24 + (h_cnt - 600)];
                end
                else begin
                    background = 1;
                    vga = 12'h000;
                end
            end
            else begin
                background = 1;
                vga = 12'h000;
            end
        end
        else begin
            if(h_cnt >= 600 && h_cnt <= 623 && v_cnt >= 10 && v_cnt <= 39) begin
                if(pause2[(v_cnt - 10) * 24 + (h_cnt - 600)] != 12'hAEF) begin
                    background = 0;
                    vga = pause2[(v_cnt - 10) * 24 + (h_cnt - 600)];
                end
                else begin
                    background = 1;
                    vga = 12'h000;
                end
            end
            else begin
                background = 1;
                vga = 12'h000;
            end
        end

    end
endmodule
/*
module bait_home (
    input [9:0] h_cnt,
    input [9:0] v_cnt,
    output reg background, //1 for print background 0 for print fish
    output reg [11:0] vga
);

    parameter [11:0] bait_home [0:719] = {//24*30

    };

    always @(*) begin
        if(h_cnt >= 308 && h_cnt <= 331 && v_cnt >= 340 && v_cnt <= 369) begin
            if(bait_home[(v_cnt - 340) * 24 + (h_cnt - 308)] != 12'hAEF) begin
                background = 0;
                vga = bait_home[(v_cnt - 340) * 24 + (h_cnt - 308)];
            end
            else begin
                background = 1;
                vga = 12'h000;
            end
        end
        else begin
            background = 1;
            vga = 12'h000;
        end
    end
endmodule*/