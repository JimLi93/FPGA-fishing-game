module shark (
    input [9:0] h_cnt,
    input [9:0] v_cnt,
    input [9:0] fish_h_position,
    input [9:0] fish_v_position,
    input fish_way,  //0 for go left , 1 for go right , 2 for go up
    input fish_appear, //1 for fish appear 0 for the fish doesn't exist
    output reg background, //1 for print background 0 for print fish
    output reg [11:0] vga
);
    parameter [11:0] shark [0:7551] = {//118*64
        //get rid of up1 line && down 1 line
        //get rid of 353,351,452,453, 463, 464 etc.
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h332,12'h232,12'h232,12'h343,12'h343,12'h343,12'h232,12'h232,12'h232,12'h343,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h332,12'h232,12'h232,12'h232,12'h232,12'h232,12'h232,12'h232,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h333,12'h233,12'h233,12'h344,12'h445,12'h445,12'h556,12'h556,12'h567,12'h567,12'h567,12'h556,12'h556,12'h556,12'h445,12'h345,12'h334,12'h233,12'h233,12'h232,12'h343,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h332,12'h333,12'h233,12'h344,12'h455,12'h566,12'h667,12'h678,12'h778,12'h778,12'h678,12'h667,12'h667,12'h556,12'h334,12'h223,12'h333,12'h332,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h233,12'h333,12'h445,12'h556,12'h668,12'h678,12'h678,12'h668,12'h668,12'h668,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h567,12'h668,12'h668,12'h678,12'h668,12'h667,12'h556,12'h445,12'h334,12'h333,12'h232,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h332,12'h233,12'h444,12'h667,12'h789,12'h889,12'h889,12'h789,12'h778,12'h678,12'h678,12'h678,12'h678,12'h678,12'h678,12'h678,12'h779,12'h778,12'h668,12'h555,12'h222,12'h110,12'h131,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h233,12'h333,12'h455,12'h667,12'h678,12'h668,12'h667,12'h667,12'h567,12'h667,12'h667,12'h667,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h667,12'h556,12'h445,12'h233,12'h233,12'h343,12'h352,12'h352,12'h352,12'h352,12'h343,12'h232,12'h334,12'h667,12'h889,12'h789,12'h678,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h567,12'h667,12'h668,12'h668,12'h667,12'h667,12'h555,12'h333,12'h232,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h232,12'h334,12'h556,12'h668,12'h668,12'h667,12'h667,12'h668,12'h667,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h668,12'h567,12'h344,12'h233,12'h333,12'h343,12'h232,12'h444,12'h667,12'h789,12'h678,12'h568,12'h567,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h667,12'h668,12'h667,12'h667,12'h667,12'h345,12'h233,12'h333,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h233,12'h334,12'h567,12'h668,12'h667,12'h667,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h567,12'h667,12'h667,12'h667,12'h667,12'h668,12'h556,12'h223,12'h223,12'h556,12'h678,12'h567,12'h668,12'h568,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h668,12'h667,12'h344,12'h232,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h233,12'h556,12'h668,12'h667,12'h668,12'h668,12'h667,12'h668,12'h667,12'h567,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h667,12'h567,12'h667,12'h667,12'h668,12'h668,12'h668,12'h668,12'h567,12'h334,12'h233,12'h556,12'h678,12'h667,12'h667,12'h667,12'h667,12'h567,12'h567,12'h667,12'h668,12'h667,12'h445,12'h232,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h233,12'h456,12'h668,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h667,12'h667,12'h678,12'h678,12'h556,12'h233,12'h334,12'h667,12'h667,12'h667,12'h567,12'h667,12'h667,12'h667,12'h556,12'h233,12'h332,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h232,12'h233,12'h455,12'h667,12'h667,12'h567,12'h667,12'h668,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h667,12'h667,12'h667,12'h567,12'h456,12'h456,12'h445,12'h445,12'h456,12'h456,12'h557,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h667,12'h667,12'h667,12'h668,12'h667,12'h678,12'h556,12'h223,12'h445,12'h678,12'h667,12'h667,12'h668,12'h444,12'h232,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h232,12'h222,12'h333,12'h444,12'h333,12'h233,12'h233,12'h233,12'h333,12'h233,12'h233,12'h344,12'h556,12'h667,12'h667,12'h667,12'h667,12'h567,12'h667,12'h567,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h568,12'h567,12'h567,12'h668,12'h779,12'h9AB,12'hBBC,12'h789,12'h667,12'h667,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h334,12'h334,12'h667,12'h667,12'h333,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h232,12'h352,12'h343,12'h232,12'h343,12'h352,
        12'h352,12'h352,12'h343,12'h233,12'h556,12'h668,12'h668,12'h668,12'h678,12'h668,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h668,12'h668,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h567,12'h789,12'hABC,12'hBCD,12'h9AB,12'h789,12'h668,12'h567,12'h667,12'h667,12'h678,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h667,12'h667,12'h567,12'h667,12'h667,12'h445,12'h223,12'h223,12'h454,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h332,12'h232,12'h445,12'h556,12'h567,12'h667,12'h556,12'h444,12'h222,
        12'h352,12'h454,12'h233,12'h667,12'h668,12'h568,12'h668,12'h668,12'h668,12'h668,12'h668,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h667,12'h667,12'h667,12'h567,12'h567,12'h668,12'h89A,12'hABC,12'h9AB,12'h789,12'h568,12'h567,12'h567,12'h678,12'h667,12'h556,12'h445,12'h334,12'h334,12'h446,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h667,12'h677,12'h567,12'h333,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h232,12'h455,12'h667,12'h667,12'h667,12'h668,12'h668,12'h667,12'h677,12'h333,
        12'h352,12'h233,12'h567,12'h668,12'h668,12'h567,12'h567,12'h567,12'h667,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h667,12'h567,12'h678,12'h99B,12'hABC,12'h89A,12'h678,12'h567,12'h567,12'h667,12'h678,12'h567,12'h344,12'h333,12'h444,12'h223,12'h556,12'h556,12'h334,12'h334,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h567,12'h667,12'h668,12'h667,12'h233,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h233,12'h567,12'h668,12'h667,12'h667,12'h667,12'h667,12'h668,12'h667,12'h556,12'h233,
        12'h352,12'h333,12'h678,12'h668,12'h789,12'h789,12'h778,12'h678,12'h567,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h678,12'h667,12'h667,12'h789,12'h89A,12'h667,12'h567,12'h567,12'h668,12'h667,12'h556,12'h334,12'h333,12'h222,12'hCCC,12'hCCC,12'h444,12'h668,12'h668,12'h668,12'h567,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h567,12'h667,12'h668,12'h667,12'h334,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h233,12'h667,12'h677,12'h667,12'h668,12'h667,12'h667,12'h667,12'h568,12'h678,12'h334,12'h454,
        12'h343,12'h445,12'h668,12'h567,12'h678,12'h88A,12'h88A,12'h789,12'h789,12'h678,12'h668,12'h567,12'h567,12'h567,12'h667,12'h667,12'h667,12'h668,12'h668,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h667,12'h678,12'h345,12'h445,12'h667,12'h567,12'h567,12'h667,12'h668,12'h667,12'h555,12'h333,12'h433,12'h433,12'h211,12'h333,12'hFEE,12'hAAA,12'h445,12'h678,12'h668,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h667,12'h667,12'h668,12'h334,12'h332,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h232,12'h567,12'h668,12'h667,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h566,12'h233,12'h352,
        12'h454,12'h445,12'h668,12'h667,12'h567,12'h678,12'h889,12'h889,12'h889,12'h88A,12'h789,12'h789,12'h678,12'h678,12'h667,12'h567,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h567,12'h667,12'h667,12'h668,12'h446,12'h234,12'h667,12'h667,12'h668,12'h678,12'h667,12'h555,12'h333,12'h322,12'h322,12'h211,12'h211,12'h101,12'h766,12'hFFF,12'h888,12'h445,12'h668,12'h667,12'h567,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h344,12'h232,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h233,12'h455,12'h668,12'h567,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h668,12'h444,12'h443,12'h352,
        12'h352,12'h445,12'h667,12'h567,12'h567,12'h567,12'h668,12'h789,12'h889,12'h789,12'h789,12'h889,12'h889,12'h889,12'h789,12'h789,12'h779,12'h678,12'h678,12'h668,12'h667,12'h667,12'h667,12'h667,12'h668,12'h567,12'h567,12'h667,12'h567,12'h223,12'h667,12'h668,12'h678,12'h667,12'h445,12'h223,12'h211,12'h211,12'h211,12'h211,12'h211,12'h211,12'h111,12'hCCC,12'hFFF,12'h556,12'h556,12'h668,12'h667,12'h567,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h568,12'h668,12'h667,12'h445,12'h333,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h334,12'h667,12'h668,12'h567,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h567,12'h233,12'h352,12'h352,
        12'h352,12'h445,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h678,12'h789,12'h88A,12'h889,12'h889,12'h789,12'h889,12'h889,12'h889,12'h789,12'h889,12'h889,12'h789,12'h778,12'h667,12'h567,12'h668,12'h667,12'h667,12'h667,12'h334,12'h666,12'h668,12'h567,12'h344,12'h334,12'h444,12'h100,12'h111,12'h211,12'h211,12'h211,12'h211,12'h110,12'h666,12'hFFF,12'hEEE,12'h334,12'h667,12'h668,12'h667,12'h567,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h568,12'h668,12'h667,12'h668,12'h446,12'h233,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h233,12'h667,12'h667,12'h668,12'h667,12'h667,12'h667,12'h667,12'h567,12'h668,12'h668,12'h445,12'h343,12'h352,12'h352,
        12'h352,12'h344,12'h678,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h567,12'h678,12'h779,12'h789,12'h889,12'h889,12'h889,12'h789,12'h889,12'h889,12'h889,12'h889,12'h88A,12'h668,12'h668,12'h668,12'h667,12'h667,12'h667,12'h223,12'h444,12'h333,12'h223,12'h555,12'hDDD,12'hEEE,12'h999,12'h444,12'h211,12'h100,12'h100,12'h111,12'h555,12'hEED,12'hFFF,12'hAAA,12'h444,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h668,12'h667,12'h668,12'h556,12'h232,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h455,12'h678,12'h667,12'h668,12'h667,12'h667,12'h667,12'h667,12'h668,12'h667,12'h667,12'h233,12'h352,12'h352,12'h352,
        12'h352,12'h233,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h567,12'h667,12'h678,12'h779,12'h789,12'h889,12'h789,12'h789,12'h889,12'h889,12'h789,12'h668,12'h668,12'h668,12'h667,12'h667,12'h667,12'h556,12'h556,12'h667,12'h667,12'h334,12'h889,12'hFFF,12'hFFF,12'hEEE,12'hCCC,12'hA99,12'h999,12'hCCC,12'hFFF,12'hFFF,12'hDDD,12'h334,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h668,12'h667,12'h668,12'h668,12'h556,12'h233,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h233,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h667,12'h455,12'h343,12'h352,12'h352,12'h352,
        12'h352,12'h233,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h567,12'h667,12'h668,12'h678,12'h678,12'h678,12'h668,12'h567,12'h668,12'h567,12'h668,12'h667,12'h667,12'h667,12'h668,12'h668,12'h668,12'h668,12'h667,12'h334,12'h778,12'hEDD,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hDDE,12'h555,12'h455,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h677,12'h566,12'h667,12'h667,12'h667,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h667,12'h667,12'h233,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h445,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h678,12'h333,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h343,12'h556,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h667,12'h667,12'h667,12'h668,12'h668,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h668,12'h568,12'h568,12'h667,12'h667,12'h445,12'h444,12'h888,12'hCCC,12'hDDD,12'hDDD,12'hCCC,12'h889,12'h444,12'h445,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h334,12'h667,12'h445,12'h556,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h667,12'h667,12'h668,12'h345,12'h333,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h233,12'h667,12'h667,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h677,12'h567,12'h333,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h343,12'h445,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h678,12'h567,12'h344,12'h233,12'h223,12'h233,12'h223,12'h444,12'h567,12'h667,12'h567,12'h667,12'h667,12'h567,12'h567,12'h567,12'h567,12'h667,12'h667,12'h667,12'h667,12'h445,12'h567,12'h445,12'h345,12'h567,12'h667,12'h668,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h678,12'h456,12'h233,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h242,12'h445,12'h667,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h445,12'h343,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h233,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h678,12'h678,12'h667,12'h677,12'h667,12'h667,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h667,12'h667,12'h456,12'h667,12'h667,12'h668,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h567,12'h668,12'h667,12'h344,12'h232,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h232,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h678,12'h334,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h233,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h668,12'h668,12'h668,12'h667,12'h567,12'h668,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h334,12'h233,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h445,12'h668,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h333,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h455,12'h668,12'h667,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h667,12'h667,12'h667,12'h667,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h667,12'h667,12'h445,12'h233,12'h233,12'h343,12'h343,12'h352,12'h352,12'h343,12'h343,12'h334,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h668,12'h445,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h334,12'h667,12'h668,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h678,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h668,12'h445,12'h556,12'h667,12'h667,12'h667,12'h668,12'h667,12'h667,12'h667,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h667,12'h668,12'h667,12'h567,12'h445,12'h334,12'h333,12'h333,12'h333,12'h455,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h668,12'h334,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h232,12'h567,12'h668,12'h667,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h677,12'h567,12'h344,12'h445,12'h334,12'h233,12'h223,12'h223,12'h333,12'h334,12'h445,12'h556,12'h667,12'h668,12'h668,12'h667,12'h567,12'h567,12'h335,12'h678,12'h667,12'h667,12'h667,12'h667,12'h567,12'h345,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h568,12'h667,12'h677,12'h667,12'h667,12'h678,12'h667,12'h667,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h567,12'h667,12'h233,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h445,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h445,12'h556,12'hCCC,12'hEEE,12'h999,12'hCCC,12'hEEE,12'hDDD,12'hCCC,12'hBBB,12'h888,12'h556,12'h334,12'h334,12'h445,12'h567,12'h667,12'h678,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h445,12'h556,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h667,12'h667,12'h232,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h233,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h668,12'h667,12'h667,12'h566,12'h233,12'h999,12'hFFF,12'hFFF,12'hFFF,12'h888,12'hDDD,12'hEEE,12'hEEE,12'hEEE,12'hEEF,12'hEEF,12'hEEF,12'hEEE,12'hCCC,12'h888,12'h344,12'h223,12'h445,12'h556,12'h334,12'h667,12'h667,12'h667,12'h667,12'h667,12'h122,12'h556,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h667,12'h667,12'h667,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h566,12'h232,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h343,12'h556,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h667,12'h667,12'h667,12'h445,12'h555,12'h667,12'h777,12'hBBB,12'hFFF,12'hFFF,12'h988,12'hDDD,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hEEE,12'hEEF,12'hEEE,12'hCCC,12'h888,12'h344,12'h334,12'h667,12'h667,12'h668,12'h667,12'h667,12'h233,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h556,12'h344,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h233,12'h667,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h567,12'h567,12'h667,12'h678,12'h567,12'h334,12'h888,12'hDDD,12'h888,12'hEEE,12'h778,12'hAAA,12'hFFF,12'h999,12'hDDD,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEF,12'hCCC,12'h334,12'h557,12'h667,12'h668,12'h667,12'h667,12'h334,12'h456,12'h668,12'h667,12'h667,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h456,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h233,12'h556,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h567,12'h567,12'h567,12'h668,12'h668,12'h667,12'h445,12'h334,12'h999,12'hFFF,12'hCCC,12'h999,12'hEEE,12'hEEE,12'h999,12'h999,12'h888,12'hDDD,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hCCC,12'h334,12'h557,12'h667,12'h667,12'h667,12'h667,12'h567,12'h223,12'h567,12'h668,12'h567,12'h668,12'h668,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h556,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h233,12'h667,12'h667,12'h568,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h667,12'h445,12'h555,12'hBBB,12'hAA9,12'h655,12'hEDD,12'h998,12'hCCC,12'hEEE,12'hDEE,12'hEEF,12'hAAB,12'h445,12'hDDD,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hBCC,12'h344,12'h556,12'h667,12'h667,12'h667,12'h668,12'h668,12'h556,12'h223,12'h567,12'h668,12'h667,12'h567,12'h567,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h567,12'h667,12'h667,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h668,12'h456,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h445,12'h668,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h668,12'h567,12'h668,12'h668,12'h668,12'h667,12'h445,12'h555,12'hAAB,12'hFFF,12'hFFF,12'h888,12'hAAA,12'h888,12'h888,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hEEF,12'hCCD,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hBCC,12'h344,12'h556,12'h667,12'h667,12'h667,12'h667,12'h668,12'h667,12'h556,12'h223,12'h444,12'h667,12'h678,12'h668,12'h668,12'h668,12'h667,12'h667,12'h567,12'h667,12'h567,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h668,12'h667,12'h567,12'h667,12'h667,12'h567,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h456,12'h344,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h232,12'h556,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h667,12'h667,12'h668,12'h667,12'h567,12'h556,12'h556,12'h667,12'h668,12'h556,12'h334,12'h556,12'h555,12'h888,12'hFEE,12'hFFF,12'hFFF,12'h777,12'hEEE,12'h999,12'h888,12'hEEF,12'hDEE,12'hEEE,12'hDDE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hBCC,12'h345,12'h556,12'h667,12'h567,12'h667,12'h667,12'h567,12'h667,12'h667,12'h566,12'h222,12'h223,12'h334,12'h445,12'h667,12'h678,12'h668,12'h668,12'h668,12'h667,12'h567,12'h567,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h567,12'h668,12'h668,12'h667,12'h668,12'h678,12'h678,12'h667,12'h667,12'h667,12'h678,12'h678,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h567,12'h556,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h233,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h557,12'h456,12'h445,12'h556,12'h667,12'h677,12'h556,12'h223,12'h344,12'hAAB,12'hEEE,12'h877,12'h999,12'h777,12'hEEE,12'hFFF,12'h777,12'hEEE,12'hEEE,12'hDDE,12'hEEE,12'hEEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hDDE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hCCC,12'h345,12'h556,12'h667,12'h567,12'h667,12'h667,12'h668,12'h567,12'h668,12'h667,12'h667,12'h333,12'hAAB,12'h666,12'h222,12'h223,12'h556,12'h678,12'h678,12'h668,12'h667,12'h567,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h678,12'h678,12'h667,12'h556,12'h334,12'h122,12'h222,12'h222,12'h222,12'h223,12'h223,12'h233,12'h567,12'h667,12'h567,12'h667,12'h667,12'h667,12'h667,12'h567,12'h667,12'h567,12'h232,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h233,12'h445,12'h677,12'h667,12'h456,12'h556,12'h556,12'h556,12'h556,12'h567,12'h667,12'h556,12'h334,12'h333,12'h555,12'h333,12'hCCC,12'hFFF,12'hEEE,12'h777,12'hEEE,12'h999,12'h888,12'hBBB,12'h999,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hCCC,12'h344,12'h556,12'h667,12'h567,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h678,12'h555,12'h556,12'hDDD,12'hCCC,12'h777,12'h444,12'h333,12'h334,12'h455,12'h556,12'h667,12'h677,12'h667,12'h667,12'h668,12'h668,12'h678,12'h678,12'h678,12'h678,12'h567,12'h556,12'h445,12'h334,12'h334,12'h445,12'h777,12'h999,12'hBBB,12'hCCC,12'hAAA,12'h222,12'h232,12'h333,12'h445,12'h678,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h667,12'h233,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h232,12'h445,12'h566,12'h556,12'h556,12'h445,12'h334,12'h223,12'h223,12'h222,12'h334,12'h999,12'hDCC,12'hBBB,12'h888,12'h777,12'hEEE,12'hCCC,12'h999,12'hEEE,12'hEEE,12'hCCD,12'h899,12'hDDD,12'hEEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hCCC,12'h334,12'h556,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h678,12'h334,12'h889,12'hEEE,12'hEEF,12'hEEE,12'hCDD,12'hAAA,12'h777,12'h445,12'h333,12'h333,12'h334,12'h334,12'h334,12'h334,12'h334,12'h333,12'h334,12'h334,12'h334,12'h555,12'h888,12'hABB,12'hDDE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hCCC,12'h444,12'h352,12'h352,12'h352,12'h333,12'h678,12'h668,12'h667,12'h667,12'h667,12'h667,12'h668,12'h567,12'h667,12'h233,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h221,12'h445,12'h667,12'h444,12'h888,12'h888,12'h999,12'hBBB,12'h877,12'h777,12'hEDD,12'hFFF,12'h777,12'hDDD,12'hAAB,12'h888,12'h888,12'hDDD,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDDD,12'h333,12'h556,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h334,12'hDDE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hFEF,12'hEEF,12'hEEE,12'hDDD,12'hBBB,12'hAAA,12'hAAA,12'h9AA,12'h9AA,12'hABB,12'hCCC,12'hDDD,12'hEEE,12'hEFF,12'hEEF,12'hEEE,12'hDEE,12'hDEE,12'hEEE,12'hEEE,12'hDDD,12'h444,12'h352,12'h352,12'h352,12'h352,12'h233,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h344,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h454,12'hDCC,12'hCCC,12'h777,12'hCCC,12'hFFF,12'hEEE,12'h888,12'hBBB,12'h999,12'hAAA,12'hAAA,12'hEEE,12'hEEF,12'h999,12'h777,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hDEE,12'hEEE,12'hEEE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hEEE,12'h334,12'h567,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h445,12'h99A,12'hEEF,12'hDEE,12'hEEE,12'hEEE,12'hDEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hEEE,12'hDEE,12'h555,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h445,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h556,12'h242,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h443,12'hDDD,12'hDDD,12'h777,12'h999,12'h989,12'hBBB,12'hEEE,12'h777,12'h777,12'hEEE,12'hDEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'h444,12'h667,12'h556,12'h668,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h567,12'h555,12'hEEF,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hEEE,12'hDEE,12'hEEE,12'hEEE,12'hEEE,12'hDEE,12'hEEE,12'hEEE,12'h677,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h344,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h233,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'hCCC,12'hFFF,12'hAAA,12'h778,12'hEEE,12'hEEE,12'hDDD,12'hDDD,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEFF,12'h555,12'h667,12'h455,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h333,12'hDDD,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hEEE,12'hDEE,12'hEEE,12'hDEE,12'hEEE,12'hEEE,12'h777,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h333,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h678,12'h344,12'h343,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h454,12'hBBB,12'hEEE,12'hEEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'h778,12'h556,12'h556,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h678,12'h344,12'hBBB,12'hEEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hEEE,12'hDEE,12'hEEE,12'hEEF,12'hDDD,12'h666,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h455,12'h667,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h556,12'h333,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h999,12'hEEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hBBB,12'h344,12'h667,12'h456,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h556,12'h777,12'hEEF,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hEEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hEEE,12'hDEE,12'hEEE,12'hEEE,12'hCCC,12'h454,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h333,12'h668,12'h667,12'h667,12'h668,12'h667,12'h667,12'h567,12'h667,12'h667,12'h233,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h443,12'h777,12'hDDD,12'hEEE,12'hEEE,12'hEEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDDE,12'h334,12'h667,12'h446,12'h667,12'h667,12'h667,12'h667,12'h567,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h445,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hEEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hEEE,12'hEEE,12'h999,12'h333,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h332,12'h455,12'h677,12'h667,12'h668,12'h667,12'h667,12'h667,12'h667,12'h668,12'h344,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h454,12'h443,12'hBBB,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hEEE,12'hEEF,12'h677,12'h556,12'h567,12'h556,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h668,12'h677,12'h223,12'hCDD,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hEEE,12'hCCC,12'h555,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h232,12'h677,12'h667,12'h668,12'h667,12'h667,12'h667,12'h667,12'h668,12'h566,12'h232,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h776,12'hDDD,12'hEEE,12'hDEE,12'h778,12'hBBB,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hCCC,12'h333,12'h667,12'h446,12'h667,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h667,12'h667,12'h344,12'hAAA,12'hEEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hEEF,12'hDEE,12'h888,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h445,12'h678,12'h568,12'h567,12'h567,12'h667,12'h567,12'h668,12'h667,12'h233,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h999,12'hEEE,12'hEEE,12'h999,12'h9AA,12'hEEE,12'hEEE,12'hEEE,12'hEEF,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hEEF,12'h667,12'h555,12'h556,12'h556,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h567,12'h667,12'h556,12'h666,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hEEE,12'hEEF,12'hBBB,12'h454,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h333,12'h556,12'h668,12'h568,12'h567,12'h667,12'h667,12'h568,12'h678,12'h344,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h454,12'hAAA,12'hEEE,12'hEEF,12'hEEE,12'hEEE,12'h999,12'hAAA,12'hDDD,12'hEEE,12'hEEF,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hEEE,12'hDDD,12'h334,12'h667,12'h456,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h677,12'h334,12'hDDE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hEEE,12'hEEF,12'hCCC,12'h555,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h233,12'h556,12'h678,12'h667,12'h668,12'h667,12'h568,12'h667,12'h556,12'h232,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h221,12'h444,12'h999,12'hEEE,12'hFEF,12'hDDD,12'hAAA,12'h777,12'h677,12'h999,12'hCCC,12'hEEE,12'hEEF,12'hEEF,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hAAB,12'h233,12'h556,12'h456,12'h668,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h677,12'h334,12'hAAB,12'hEEE,12'hEEE,12'hDEE,12'hEEE,12'hEEE,12'hEEE,12'hBBC,12'h566,12'h332,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h233,12'h334,12'h566,12'h678,12'h667,12'h668,12'h668,12'h667,12'h233,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h444,12'h667,12'h344,12'h334,12'h778,12'hCCC,12'hFFF,12'hFFF,12'hDDE,12'hBBB,12'h889,12'h777,12'h778,12'hAAA,12'hCCC,12'hDDE,12'hEEF,12'hEEF,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hDEE,12'hEEE,12'hEEE,12'hEEE,12'hDEE,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hEEE,12'h888,12'h334,12'h556,12'h667,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h566,12'h556,12'hEEE,12'hEEE,12'hEEF,12'hDDE,12'hAAA,12'h565,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h233,12'h333,12'h444,12'h556,12'h567,12'h667,12'h344,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h455,12'h667,12'h668,12'h667,12'h455,12'h334,12'h445,12'h888,12'hCCC,12'hEEF,12'hFFF,12'hEEF,12'hDDD,12'hBBB,12'h999,12'h777,12'h667,12'h778,12'h999,12'hAAB,12'hBBC,12'hCCD,12'hDDD,12'hDDE,12'hDDE,12'hDDD,12'hDDD,12'hCCC,12'hDDE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hDEE,12'hEEE,12'h778,12'h334,12'h455,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h334,12'hBBB,12'hBBB,12'h777,12'h444,12'h454,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h232,12'h333,12'h222,12'h242,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h232,12'h455,12'h667,12'h668,12'h667,12'h668,12'h678,12'h334,12'h232,12'h343,12'h555,12'h888,12'hBBB,12'hDDD,12'hEFF,12'hFFF,12'hFFF,12'hEEE,12'hCCD,12'hBBB,12'hAAA,12'h999,12'h888,12'h888,12'h888,12'h878,12'h778,12'h788,12'h888,12'hCCD,12'hEEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hDEE,12'hEEE,12'hEEE,12'h667,12'h334,12'h456,12'h668,12'h667,12'h667,12'h667,12'h667,12'h667,12'h667,12'h668,12'h456,12'h333,12'h443,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h232,12'h556,12'h667,12'h668,12'h667,12'h678,12'h445,12'h343,12'h352,12'h352,12'h352,12'h343,12'h343,12'h444,12'h555,12'h777,12'h9AA,12'hBBB,12'hDDD,12'hEEF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFFF,12'hFEF,12'hEEE,12'hEEE,12'hEEF,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'h666,12'h333,12'h556,12'h667,12'h568,12'h568,12'h667,12'h667,12'h667,12'h667,12'h667,12'h334,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h567,12'h667,12'h667,12'h678,12'h445,12'h232,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h343,12'h352,12'h444,12'h555,12'h777,12'h888,12'h999,12'h99A,12'hBAB,12'hBBC,12'hCCC,12'hCCC,12'hDDD,12'hDDD,12'hCDD,12'hCCC,12'hCCC,12'hCCC,12'hBBB,12'hAAA,12'h999,12'h888,12'h777,12'h555,12'h221,12'h222,12'h556,12'h678,12'h667,12'h667,12'h667,12'h668,12'h667,12'h667,12'h556,12'h233,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h567,12'h668,12'h668,12'h445,12'h231,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h564,12'h232,12'h352,12'h443,12'h564,12'h565,12'h676,12'h676,12'h675,12'h665,12'h565,12'h454,12'h352,12'h332,12'h332,12'h564,12'h352,12'h352,12'h352,12'h232,12'h112,12'h556,12'h667,12'h667,12'h667,12'h668,12'h668,12'h567,12'h667,12'h334,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h454,12'h667,12'h678,12'h445,12'h232,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h222,12'h445,12'h667,12'h667,12'h567,12'h567,12'h668,12'h667,12'h567,12'h233,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h454,12'h678,12'h445,12'h232,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h232,12'h334,12'h667,12'h668,12'h667,12'h668,12'h567,12'h678,12'h455,12'h232,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h333,12'h344,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h233,12'h445,12'h667,12'h668,12'h668,12'h668,12'h667,12'h344,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h121,12'h232,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h233,12'h446,12'h667,12'h678,12'h667,12'h667,12'h233,12'h454,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h232,12'h344,12'h455,12'h667,12'h667,12'h333,12'h443,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h233,12'h232,12'h333,12'h444,12'h221,12'h232,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h232,12'h121,12'h241,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352

    };


    always @(*) begin
        if(fish_appear == 1'b0) begin
            background = 1;
            vga = 12'h000;
        end
        else if(fish_way == 0) begin
            if(((h_cnt + 118) - fish_h_position) <= 117 && (v_cnt - fish_v_position) <= 63) begin
                if(shark[(v_cnt - fish_v_position) * 118 + (h_cnt + 118 - fish_h_position)] != 12'h352) begin
                    background = 0;
                    vga = shark[(v_cnt - fish_v_position) * 118 + (h_cnt + 118 - fish_h_position)];
                end
                else begin
                    background = 1;
                    vga = 12'h000;
                end
            end
            else begin
                background = 1;
                vga = 12'h000;
            end
        end
        else if(fish_way == 1) begin
            if(((h_cnt + 118) - fish_h_position) <= 117 && (v_cnt - fish_v_position) <= 63) begin
                if(shark[(v_cnt - fish_v_position) * 118 + (fish_h_position - h_cnt - 1)] != 12'h352) begin
                    background = 0;
                    vga = shark[(v_cnt - fish_v_position) * 118 + (fish_h_position - h_cnt - 1)];
                end
                else begin
                    background = 1;
                    vga = 12'h000;
                end
            end
            else begin
                background = 1;
                vga = 12'h000;
            end
        end
        else begin
            background = 1;
            vga = 12'h000;
        end

    end
    
endmodule

module mouth (
    input [9:0] h_cnt,
    input [9:0] v_cnt,
    input [2:0] type,
    output reg background, //1 for print background 0 for print fish
    output reg [11:0] vga
);
    parameter [11:0] mouth [0:2719] = {//40*68
        //get rid of up1 line && down 1 line
        //get rid of 353,351,452,453, 463, 464 etc.
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h111,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h222,12'h777,12'h555,12'h111,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h333,12'h888,12'h999,12'h999,12'h666,12'h111,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h444,12'h888,12'hA99,12'hCCC,12'hBBB,12'h999,12'h777,12'h111,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h333,12'h888,12'hAAA,12'hEEE,12'hEEE,12'hEEE,12'hCCC,12'h999,12'h666,12'h111,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h222,12'h888,12'hA99,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hBBB,12'h999,12'h666,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h111,12'h777,12'h999,12'hDDD,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hAAA,12'h888,12'h444,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h555,12'h999,12'hBBB,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hDDD,12'h999,12'h888,12'h222,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h222,12'h888,12'h999,12'hEED,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hAAA,12'h999,12'h666,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h666,12'h999,12'hBBB,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hDDD,12'h999,12'h888,12'h333,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h333,12'h888,12'h999,12'hEDD,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hAAA,12'h999,12'h666,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h666,12'h999,12'hAAA,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hDDC,12'h999,12'h888,12'h333,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h222,12'h777,12'h999,12'hDCC,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'h999,12'h999,12'h555,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h444,12'h888,12'h999,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hBBB,12'h999,12'h777,12'h111,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h666,12'h999,12'hBBB,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hDDD,12'h999,12'h888,12'h333,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h111,12'h777,12'h999,12'hDDD,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'h999,12'h999,12'h555,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h222,12'h888,12'h999,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hBBB,12'h999,12'h777,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h333,12'h888,12'hBAA,12'hEEE,12'hEEE,12'hEEE,12'hFEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hFEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hDCC,12'h999,12'h888,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h222,12'h444,12'h989,12'hCCC,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hCDD,12'hBCC,12'hACC,12'hACC,12'hBCD,12'hDDD,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'h999,12'h888,12'h333,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h111,12'h878,12'h555,12'h999,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hDDD,12'hDDD,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hDEE,12'hCDD,12'hDEE,12'hEEE,12'hEEE,12'hFEE,12'hAAA,12'h988,12'h666,12'h666,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h222,12'h666,12'h888,12'hAAA,12'hFEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hDDD,12'hDDD,12'hDDD,12'hDDD,12'hDDD,12'hDDD,12'hEEE,12'hEEE,12'hEEE,12'hFEE,12'hEEE,12'hCCC,12'h999,12'h888,12'h222,12'h222,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h222,12'h000,12'h444,12'h999,12'hBBB,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hDDD,12'h999,12'h888,12'h000,12'h222,12'h111,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h444,12'hAAA,12'h555,12'h777,12'hDDD,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hCCC,12'h9AA,12'h9AA,12'hAAA,12'hBBB,12'hDDD,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'h999,12'h777,12'h222,12'h777,12'h444,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h222,12'h333,12'h000,12'h777,12'h555,12'hEEE,12'hEEE,12'hEEE,12'hEEE,12'hCDD,12'h666,12'h311,12'h401,12'h611,12'h611,12'h511,12'h501,12'h311,12'h444,12'h9AA,12'hEEE,12'hEEE,12'hEEE,12'hFEE,12'h999,12'h666,12'h333,12'h222,12'h666,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h444,12'h444,12'h444,12'h988,12'h666,12'hEEE,12'hEEE,12'hEEE,12'h899,12'h311,12'h811,12'hA11,12'hA22,12'hA22,12'hA11,12'hA11,12'hA22,12'hA11,12'h911,12'h511,12'h444,12'hCDD,12'hEEE,12'hEEE,12'hBBB,12'h555,12'h777,12'h111,12'h888,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h555,12'h999,12'h999,12'h777,12'hA99,12'hEEE,12'hEEE,12'h677,12'h511,12'hA22,12'hA22,12'hB77,12'hBBB,12'hBAA,12'hB22,12'hB66,12'hBBB,12'hBAA,12'hA33,12'hA23,12'h911,12'h322,12'hBCC,12'hEEE,12'hDCC,12'h555,12'h999,12'h999,12'h999,12'h111,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h555,12'h999,12'h999,12'h888,12'hDCC,12'hEEE,12'h778,12'h611,12'hA55,12'hBBA,12'hB88,12'hDBB,12'hFFF,12'hBAA,12'h933,12'h955,12'hBBB,12'hDDD,12'hB55,12'hBBB,12'hB88,12'h922,12'h322,12'hCCD,12'hEED,12'h888,12'h888,12'h999,12'h999,12'h111,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h555,12'h999,12'h999,12'h999,12'hEED,12'hABB,12'h411,12'hA11,12'hBAA,12'hDDD,12'hB99,12'h844,12'hFFF,12'hA77,12'h611,12'h611,12'hDCC,12'hDBB,12'hA44,12'hDDD,12'hEEE,12'hA55,12'h911,12'h444,12'hEEE,12'hA99,12'h999,12'h999,12'h999,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h444,12'h999,12'h999,12'h999,12'hDEE,12'h433,12'hA22,12'hB66,12'hC77,12'hFFF,12'hB99,12'h611,12'hA77,12'h822,12'h811,12'h811,12'hA66,12'h832,12'h722,12'hFFF,12'hEDD,12'hA33,12'hB55,12'h611,12'h999,12'hCBB,12'h999,12'h999,12'h989,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h444,12'h999,12'h999,12'hBAA,12'h899,12'h611,12'hCBB,12'hDCC,12'h611,12'h966,12'hA55,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'hB88,12'h722,12'hB77,12'hDDD,12'hA55,12'h433,12'hDDD,12'h999,12'h999,12'h888,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h333,12'h999,12'h999,12'hCCC,12'h433,12'hA33,12'hEEE,12'hFFF,12'h722,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'hB99,12'hFFF,12'hB88,12'h611,12'h9AA,12'hAAA,12'h999,12'h888,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h333,12'h999,12'hAAA,12'hAAB,12'h611,12'hB55,12'h955,12'hDBB,12'h933,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'hB77,12'hA88,12'hA44,12'hA33,12'h445,12'hCCB,12'h999,12'h878,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h222,12'h444,12'h999,12'hDDD,12'h555,12'hA55,12'hEEE,12'h843,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h711,12'hCAA,12'hBAA,12'h511,12'hBCC,12'h999,12'h877,12'h333,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h666,12'h888,12'hAAA,12'hDDD,12'h411,12'hB56,12'hFEE,12'hB77,12'h811,12'h811,12'h811,12'h811,12'h811,12'h711,12'h711,12'h611,12'h711,12'h711,12'h711,12'h811,12'h811,12'h811,12'h811,12'h811,12'hEEE,12'hCAA,12'h811,12'h788,12'hAAA,12'h888,12'h777,12'h222,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h111,12'h888,12'h999,12'hCCC,12'h999,12'h833,12'hBAA,12'h722,12'h822,12'h811,12'h811,12'h811,12'h611,12'h610,12'h510,12'h510,12'h510,12'h510,12'h510,12'h510,12'h610,12'h711,12'h811,12'h811,12'h811,12'h822,12'h855,12'hB88,12'h444,12'hCCC,12'h999,12'h988,12'h555,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h333,12'h999,12'h999,12'hEDD,12'h555,12'hB88,12'hFFF,12'h943,12'h811,12'h811,12'h711,12'h610,12'h510,12'h510,12'h510,12'h510,12'h610,12'h610,12'h510,12'h511,12'h610,12'h510,12'h610,12'h811,12'h811,12'h811,12'hBAA,12'hDDD,12'h423,12'hCDD,12'h999,12'h999,12'h777,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h444,12'h999,12'h999,12'hEEE,12'h422,12'hA33,12'hB77,12'h933,12'h811,12'h711,12'h510,12'h510,12'h610,12'h611,12'h711,12'h811,12'h811,12'h811,12'h811,12'h711,12'h611,12'h510,12'h510,12'h610,12'h811,12'h811,12'hA66,12'hA56,12'h711,12'hAAA,12'hAAA,12'h999,12'h888,12'h111,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h666,12'h999,12'hBAA,12'hCDC,12'h511,12'hCAA,12'h944,12'h811,12'h711,12'h510,12'h610,12'h711,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h711,12'h611,12'h610,12'h610,12'h811,12'h811,12'hBAA,12'h944,12'h777,12'hCCC,12'h999,12'h888,12'h222,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h777,12'h999,12'hBBB,12'hAAA,12'h711,12'hA55,12'hA44,12'h811,12'h611,12'h611,12'h811,12'h811,12'h811,12'h711,12'h611,12'h611,12'h610,12'h610,12'h611,12'h711,12'h711,12'h811,12'h811,12'h711,12'h610,12'h611,12'h811,12'hA66,12'hA33,12'h555,12'hEEE,12'h999,12'h999,12'h333,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h111,12'h777,12'h999,12'hCCC,12'h888,12'h944,12'hB99,12'h811,12'h711,12'h610,12'h811,12'h811,12'h711,12'h610,12'h510,12'h510,12'h510,12'h610,12'h510,12'h510,12'h510,12'h510,12'h611,12'h711,12'h811,12'h711,12'h610,12'h811,12'h833,12'hCAA,12'h533,12'hFEE,12'hA99,12'h999,12'h555,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h222,12'h888,12'h999,12'hDCC,12'h777,12'hA33,12'hA55,12'h811,12'h611,12'h811,12'h811,12'h611,12'h610,12'h611,12'h711,12'h711,12'h811,12'h811,12'h811,12'h811,12'h711,12'h711,12'h611,12'h610,12'h711,12'h811,12'h711,12'h711,12'h933,12'hB55,12'h522,12'hEEE,12'hAAA,12'h999,12'h666,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h222,12'h888,12'h999,12'hDCC,12'h666,12'hB77,12'hA66,12'h811,12'h811,12'h811,12'h711,12'h711,12'h811,12'h811,12'h811,12'h811,12'h711,12'h711,12'h711,12'h711,12'h811,12'h811,12'h811,12'h811,12'h711,12'h711,12'h811,12'h711,12'h811,12'hCBB,12'h511,12'hEEE,12'hBBB,12'h999,12'h666,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h222,12'h888,12'h999,12'hCCC,12'h655,12'hA33,12'h822,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h711,12'h610,12'h510,12'h510,12'h510,12'h510,12'h510,12'h510,12'h611,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'hA44,12'h511,12'hEEE,12'hBBB,12'h999,12'h666,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h222,12'h777,12'h999,12'hCCC,12'h666,12'hA22,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h611,12'h711,12'h711,12'h811,12'h811,12'h811,12'h811,12'h811,12'h711,12'h711,12'h611,12'h711,12'h811,12'h811,12'h811,12'h811,12'h811,12'h911,12'h511,12'hEEE,12'hBAA,12'h999,12'h666,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h111,12'h777,12'h999,12'hBBB,12'h777,12'hA22,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h711,12'h611,12'h610,12'h611,12'h610,12'h610,12'h711,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'h811,12'hA11,12'h522,12'hEEE,12'hAAA,12'h999,12'h555,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h777,12'h999,12'hAAA,12'h999,12'h822,12'hB77,12'h821,12'h811,12'h811,12'h811,12'h811,12'h711,12'h610,12'h510,12'h510,12'h510,12'h510,12'h510,12'h510,12'h510,12'h610,12'h611,12'h811,12'h811,12'h811,12'h811,12'h811,12'hA55,12'hA33,12'h544,12'hEEE,12'h999,12'h888,12'h333,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h555,12'h999,12'h999,12'hCCC,12'h511,12'hB88,12'h944,12'h811,12'h811,12'h811,12'h711,12'h510,12'h611,12'h711,12'h811,12'h811,12'h811,12'h811,12'h811,12'h711,12'h611,12'h610,12'h610,12'h811,12'h811,12'h811,12'h933,12'hA55,12'hA55,12'h777,12'hEDD,12'h999,12'h888,12'h222,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h222,12'h888,12'h999,12'hEEE,12'h533,12'hA45,12'hEDD,12'h811,12'h811,12'h811,12'h711,12'h911,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'h911,12'h811,12'h711,12'h811,12'h811,12'hB77,12'hBAA,12'h711,12'hBBB,12'hCCC,12'h999,12'h666,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h777,12'h999,12'hDDD,12'h888,12'h822,12'hA77,12'hB88,12'h811,12'h811,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'h912,12'h811,12'hA54,12'hA66,12'hB66,12'h512,12'hEEE,12'hBAA,12'h999,12'h333,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h444,12'h999,12'hCBB,12'hEDD,12'h411,12'hC77,12'hDCC,12'h811,12'h811,12'h911,12'hA11,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'h811,12'h811,12'hA66,12'hCCC,12'hA22,12'h666,12'hEEE,12'h999,12'h878,12'h000,12'h111,12'h222,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h888,12'hAAA,12'hFEE,12'h777,12'h922,12'h967,12'hDBB,12'h811,12'h811,12'h911,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'h911,12'h811,12'hB77,12'hA77,12'hB66,12'h611,12'hCCB,12'hDDD,12'h999,12'h444,12'h000,12'h666,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h444,12'h999,12'hEEE,12'hDDD,12'h411,12'hB77,12'hCCC,12'h811,12'h811,12'h811,12'h911,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'h911,12'h811,12'h811,12'hB77,12'hCBB,12'hA22,12'h544,12'hEEE,12'hCBB,12'h888,12'h000,12'h000,12'hBBB,12'h333,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h777,12'hEED,12'hEEE,12'h777,12'h822,12'h955,12'hCAA,12'hA55,12'h811,12'h811,12'h911,12'hA12,12'hA12,12'hA12,12'hA12,12'hA12,12'hA11,12'h911,12'h811,12'h811,12'hCBB,12'h955,12'hB44,12'h511,12'hBBB,12'hEEE,12'hAAA,12'h333,12'h000,12'h333,12'h444,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h222,12'hDCC,12'hEEE,12'hDDD,12'h422,12'hB66,12'hEEE,12'h966,12'hA66,12'h811,12'h811,12'h811,12'h911,12'h911,12'h911,12'h911,12'h811,12'h811,12'h822,12'h955,12'hEDD,12'hBAA,12'h811,12'h666,12'hFEE,12'hEED,12'h777,12'h000,12'h000,12'h111,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h777,12'hEEE,12'hEEE,12'h999,12'h622,12'hB99,12'h855,12'hFFF,12'h944,12'h811,12'hA66,12'hB88,12'h811,12'h822,12'hDCC,12'h811,12'h811,12'hDBB,12'hA99,12'hCAA,12'hA66,12'h322,12'hDDD,12'hEEE,12'hCCC,12'h111,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hDDD,12'hEEE,12'hEEE,12'h566,12'h711,12'hA44,12'hFFF,12'hA99,12'h611,12'hDCC,12'hFEE,12'h811,12'hA66,12'hFFF,12'hA66,12'h844,12'hFFF,12'hCAA,12'hA33,12'h300,12'h001,12'h666,12'hEED,12'h666,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h999,12'hEEE,12'hEEE,12'hDDD,12'h455,12'h711,12'hBAA,12'hBBB,12'h844,12'hEEE,12'hFFF,12'h844,12'hBAA,12'hFFF,12'hCBB,12'hB99,12'hDDD,12'hA55,12'h300,12'h000,12'h000,12'h000,12'h666,12'h222,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h322,12'hEEE,12'hEEE,12'hEEE,12'hCDD,12'h556,12'h511,12'hA44,12'hB44,12'hBBB,12'hDDD,12'hA66,12'hBAA,12'hDDD,12'hC99,12'hB44,12'h933,12'h200,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h988,12'hEEE,12'hDDD,12'h777,12'h677,12'h567,12'h301,12'h911,12'hA33,12'hB55,12'hB33,12'hA33,12'hA55,12'hA22,12'h711,12'h222,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h101,12'h888,12'h111,12'h000,12'h000,12'h566,12'h89A,12'h444,12'h311,12'h611,12'h711,12'h711,12'h611,12'h200,12'h112,12'h222,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h111,12'hCCD,12'hABC,12'h9BB,12'h788,12'h667,12'h455,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h988,12'hEEE,12'hCDD,12'hBCD,12'hACC,12'h444,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h111,12'hBBB,12'hFEE,12'hEEE,12'hEEE,12'h111,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h333,12'h111,12'h111,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,
        12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000
    };


    always @(*) begin
        if(type == 0) begin
            if(h_cnt >= 300 && h_cnt <= 339 && v_cnt >= 206 && v_cnt <= 273) begin
                background = 0;
                vga = mouth[(v_cnt - 206) * 40 + (h_cnt - 300)];
            end
            else begin
                background = 1;
                vga = 12'h000;
            end
        end
        else if(type == 1) begin
            if(h_cnt >= 280 && h_cnt <= 359 && v_cnt >= 172 && v_cnt <= 307) begin
                background = 0;
                vga = mouth[((v_cnt - 172)>>1) * 40 + ((h_cnt - 280)>>1)];
            end
            else begin
                background = 1;
                vga = 12'h000;
            end
        end
        else if(type == 2) begin
            if(h_cnt >= 260 && h_cnt <= 379 && v_cnt >= 138 && v_cnt <= 341) begin
                background = 0;
                vga = mouth[((v_cnt - 138) / 3) * 40 + ((h_cnt - 260) / 3)];
            end
            else begin
                background = 1;
                vga = 12'h000;
            end
        end
        else if(type == 3) begin
            if(h_cnt >= 240 && h_cnt <= 399 && v_cnt >= 104 && v_cnt <= 375) begin
                background = 0;
                vga = mouth[((v_cnt - 104)>>2) * 40 + ((h_cnt - 240)>>2)];
            end
            else begin
                background = 1;
                vga = 12'h000;
            end
        end
        else if(type == 4) begin
            if(h_cnt >= 220 && h_cnt <= 419 && v_cnt >= 70 && v_cnt <= 409) begin
                background = 0;
                vga = mouth[((v_cnt - 70) / 5) * 40 + ((h_cnt - 220) / 5)];
            end
            else begin
                background = 1;
                vga = 12'h000;
            end
        end
        else if(type == 5) begin
            if(h_cnt >= 200 && h_cnt <= 439 && v_cnt >= 36 && v_cnt <= 443) begin
                background = 0;
                vga = mouth[((v_cnt - 36) / 6) * 40 + ((h_cnt - 200) / 6)];
            end
            else begin
                background = 1;
                vga = 12'h000;
            end
        end
        else if(type == 6) begin
            background = 0; //all black
            vga = 12'h000;
        end
        else begin
            background = 1;
            vga = 12'h000;
        end
    end
endmodule
