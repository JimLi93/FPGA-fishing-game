module fast (
    input [9:0] h_cnt,
    input [9:0] v_cnt,
    input [9:0] fish_h_position,
    input [9:0] fish_v_position,
    input fish_way,  //0 for go left , 1 for go right , 2 for go up
    input fish_appear, //1 for fish appear 0 for the fish doesn't exist
    output reg background, //1 for print background 0 for print fish
    output reg [11:0] vga
);
    parameter [11:0] fast [0:1130] = {//39*29
        //get rid of up1 line && down 1 line
        //get rid of 353,351,452,453, 463, 464 etc.
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h320,12'h430,12'h330,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h430,12'hD83,12'hD62,12'hE52,12'hD63,12'h341,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h973,12'hE72,12'hB53,12'h721,12'hD62,12'hB53,12'h343,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h343,12'h352,12'h340,12'h352,12'h552,12'h661,12'h841,12'h942,12'hB53,12'h930,12'hC53,12'h731,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h671,12'h881,12'hDE1,12'hEE1,12'hED2,12'hED2,12'hED3,12'hEE2,12'hAB2,12'hBB1,12'h851,12'hA43,12'h432,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h551,12'hDE2,12'hED1,12'hDD1,12'h752,12'h947,12'h948,12'h948,12'hA48,12'hA49,12'h947,12'hEC2,12'hEE0,12'hCD1,12'h440,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h430,12'h530,12'h341,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h230,12'hBB2,12'hEE0,12'hED0,12'hFC0,12'hFC0,12'hEC1,12'h947,12'h949,12'h948,12'h948,12'h948,12'h948,12'h852,12'hFC0,12'hED0,12'hDE0,12'h771,12'h352,12'h352,12'h352,12'h352,12'h352,12'h641,12'hE73,12'hE62,12'hD74,12'h341,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h330,12'hDE1,12'hEE0,12'hEC0,12'hFC0,12'hFC0,12'hFC0,12'hFC0,12'h851,12'h947,12'h948,12'h948,12'h948,12'h948,12'h837,12'hEC1,12'hFC0,12'hEC0,12'hED0,12'h670,12'h352,12'h352,12'h352,12'h540,12'hE73,12'hE62,12'hD62,12'hF52,12'h631,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h340,12'hCD2,12'hDC2,12'hEC0,12'hEC0,12'hEC0,12'hFC0,12'hFC0,12'hFC0,12'hEC1,12'h847,12'h939,12'h948,12'h948,12'h948,12'h947,12'h971,12'hFC0,12'hFC0,12'hFC0,12'hDC2,12'h352,12'h352,12'h441,12'hE93,12'hE52,12'h831,12'hD64,12'hA51,12'hC63,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h341,12'hDE1,12'hC95,12'h948,12'h522,12'hDA2,12'hEC0,12'hEC0,12'hFC0,12'hFC0,12'hFC0,12'h520,12'h948,12'h948,12'h948,12'h948,12'h948,12'h733,12'hFC0,12'hEC0,12'hFC0,12'hEC1,12'hBB4,12'h352,12'h863,12'hD62,12'hD53,12'hC62,12'h720,12'hC53,12'hE53,12'h341,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'hDE2,12'hDC4,12'hA48,12'h948,12'h948,12'h948,12'h962,12'hEC0,12'hFC0,12'hFC0,12'hFC0,12'hDB3,12'h947,12'h948,12'h948,12'h948,12'h948,12'h847,12'hFC1,12'hFC0,12'hFC0,12'hFC0,12'h743,12'hDC6,12'hDB4,12'hCB7,12'h742,12'hC63,12'hB53,12'h721,12'h931,12'h331,
        12'h352,12'h352,12'h352,12'h231,12'h241,12'h352,12'h781,12'hCC3,12'h746,12'h948,12'hA49,12'h948,12'h948,12'h948,12'h972,12'hFC0,12'hFC0,12'hFC0,12'hEC1,12'h836,12'h948,12'h948,12'h948,12'h948,12'h948,12'hC91,12'hFC0,12'hFC0,12'hFC0,12'h970,12'h948,12'hA47,12'hA47,12'h948,12'h611,12'hC53,12'hC53,12'hD52,12'h420,
        12'h352,12'h242,12'hCCC,12'hDEF,12'hCDE,12'h898,12'hBCB,12'hDEE,12'hDDE,12'h99A,12'h947,12'h948,12'h948,12'h948,12'h947,12'hEB2,12'hFC0,12'hFC0,12'hEC0,12'h522,12'h948,12'h948,12'h948,12'h948,12'h948,12'h861,12'hFC0,12'hFC0,12'hFC0,12'hEC2,12'h948,12'hA48,12'h948,12'h948,12'h836,12'hB52,12'hA42,12'hC42,12'h420,
        12'h352,12'hABB,12'hDEF,12'hEEF,12'hDEE,12'hBCC,12'hDEE,12'hEEF,12'hDEE,12'hDEE,12'h556,12'h948,12'h948,12'h948,12'h948,12'h521,12'hEC0,12'hFC0,12'hFC0,12'h861,12'h948,12'hA48,12'h948,12'h948,12'h948,12'h732,12'hFC0,12'hFC0,12'hFC0,12'hEC0,12'h947,12'h948,12'h948,12'hA38,12'h836,12'hA41,12'h621,12'hC52,12'h330,
        12'h352,12'hDEE,12'hEEF,12'hFFF,12'h888,12'hDEE,12'hEEF,12'hFFF,12'hEFF,12'hDEF,12'hDDE,12'h746,12'h948,12'h948,12'h948,12'h848,12'hEC0,12'hFC0,12'hFC0,12'hDB3,12'h948,12'hA48,12'h948,12'h948,12'h948,12'h632,12'hEC0,12'hEC0,12'hEC0,12'hFC0,12'h622,12'h938,12'h927,12'hA28,12'h601,12'hD52,12'hD62,12'hE51,12'h331,
        12'h241,12'hDEF,12'h888,12'h444,12'h899,12'hDEE,12'hEEF,12'h333,12'hFFF,12'hEEF,12'hDEE,12'h524,12'hA48,12'h948,12'h948,12'h948,12'hEC1,12'hFC0,12'hFC0,12'hEC1,12'h947,12'h948,12'h948,12'h949,12'h948,12'h632,12'hFC0,12'hFC0,12'hEC0,12'hEB1,12'h520,12'hB37,12'hB28,12'h937,12'hB52,12'h832,12'h731,12'hC63,12'h352,
        12'h352,12'hDDE,12'h888,12'hDDD,12'h99A,12'hDEF,12'hFFE,12'h111,12'hFFF,12'hEFF,12'hDEE,12'h524,12'h948,12'hA48,12'hA38,12'h948,12'hEC2,12'hFC0,12'hFC0,12'hEC0,12'h847,12'hA48,12'h948,12'hA48,12'h948,12'h733,12'hEA1,12'hEA1,12'hEA1,12'hEA2,12'h971,12'hB28,12'hA37,12'h823,12'h931,12'hC53,12'hE52,12'h951,12'h352,
        12'h352,12'h676,12'hDEE,12'hDEE,12'h676,12'hDEE,12'hEEF,12'hEEF,12'hEEF,12'hDEE,12'hCDD,12'h947,12'h949,12'h948,12'hA48,12'h947,12'hEC1,12'hFC0,12'hFC0,12'hEC0,12'h735,12'h938,12'h837,12'h927,12'h838,12'h733,12'hEA1,12'hEA1,12'hEA1,12'hEA1,12'hC93,12'h936,12'h833,12'h832,12'h832,12'h843,12'h942,12'h320,12'h352,
        12'h352,12'h352,12'h787,12'hCDE,12'hCCE,12'hBBB,12'hDEF,12'hDEE,12'hDEE,12'hDEE,12'h525,12'h927,12'h928,12'h838,12'h828,12'h624,12'hEA1,12'hEA1,12'hEA1,12'hEA1,12'h624,12'h828,12'h837,12'h927,12'h828,12'h743,12'hEA1,12'hEA1,12'hEA1,12'hDA1,12'hB82,12'h533,12'h442,12'h743,12'h832,12'h932,12'h632,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h341,12'h873,12'h667,12'hDDD,12'hCCC,12'h635,12'hB27,12'h938,12'h828,12'h837,12'h827,12'h521,12'hEA1,12'hEA1,12'hEA1,12'hEA1,12'h522,12'h828,12'h837,12'h927,12'h828,12'h852,12'hEA1,12'hEA1,12'hEA1,12'hD91,12'hA83,12'h432,12'h352,12'h352,12'h421,12'h421,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h231,12'h330,12'h993,12'hEC1,12'hB82,12'hA83,12'h947,12'hA27,12'h837,12'h827,12'h828,12'h828,12'h737,12'hCA3,12'hEA1,12'hEA1,12'hEA1,12'hEA1,12'h623,12'h928,12'h828,12'h828,12'h837,12'hB72,12'hEA1,12'hEA1,12'hEA2,12'hB81,12'hA84,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h341,12'hDD2,12'hED1,12'hED1,12'hEC0,12'hEA1,12'hEA1,12'hEA2,12'h622,12'h827,12'h838,12'h838,12'h827,12'h827,12'h512,12'hEA1,12'hEA1,12'hEA1,12'hEA1,12'hDA1,12'h624,12'h828,12'h837,12'h828,12'h837,12'hD92,12'hEA1,12'hDA2,12'hB82,12'hB82,12'h320,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h341,12'hDC0,12'hEA1,12'hEA2,12'hEA2,12'hEA1,12'hA71,12'hEA0,12'h962,12'h828,12'h828,12'h828,12'h827,12'h837,12'hDA3,12'hEA1,12'hDA1,12'hEA1,12'hEA1,12'hEA2,12'h735,12'h735,12'h837,12'h837,12'h837,12'hEB2,12'hC92,12'hB82,12'hB82,12'h752,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h341,12'hCA3,12'hEA1,12'hEA1,12'hEA2,12'hB93,12'h962,12'hEA1,12'h962,12'h828,12'h837,12'h927,12'h928,12'h742,12'hEA1,12'hEA1,12'hEA1,12'hEA1,12'hEA0,12'hDA2,12'hE93,12'hE83,12'hD94,12'h953,12'h522,12'hB83,12'hA82,12'hB82,12'h642,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h331,12'h972,12'hB82,12'hA83,12'h640,12'hB82,12'hB81,12'h733,12'hA37,12'h828,12'h828,12'h624,12'hEA2,12'hEA1,12'hEA1,12'hEA1,12'hEA1,12'hEA1,12'hDA3,12'hD62,12'hC52,12'h731,12'hA43,12'hD72,12'h851,12'hB83,12'h521,12'hC52,12'h842,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h873,12'hB82,12'h751,12'h834,12'hC27,12'hB28,12'h937,12'hC93,12'hEA1,12'hEA1,12'hEA1,12'hEA1,12'hEA1,12'hDA1,12'h850,12'hD63,12'hA30,12'h931,12'hB52,12'hE52,12'hB63,12'h843,12'hB53,12'hB42,12'hE53,12'h341,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h341,12'h330,12'h352,12'h432,12'h837,12'hA35,12'hB83,12'hB82,12'hB82,12'hB82,12'hC82,12'hC82,12'hB81,12'hB82,12'h731,12'hD63,12'hB52,12'hD63,12'hD63,12'hE62,12'h731,12'hC53,12'hB41,12'hA41,12'hC53,12'h341,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h442,12'h874,12'hB83,12'hB82,12'hB82,12'hB82,12'hB82,12'hB82,12'hB82,12'hB82,12'h952,12'h832,12'hC64,12'hA42,12'hD53,12'hC63,12'h632,12'h933,12'hA43,12'h832,12'h220,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,
        12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h341,12'h220,12'h530,12'h752,12'h651,12'h430,12'h320,12'h330,12'h441,12'h341,12'h732,12'h832,12'h733,12'h221,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352,12'h352
    };


    always @(*) begin
        if(fish_appear == 1'b0) begin
            background = 1;
            vga = 12'h000;
        end
        else if(fish_way == 0) begin
            if(((h_cnt + 39) - fish_h_position) <= 38 && (v_cnt - fish_v_position) <= 28) begin
                if(fast[(v_cnt - fish_v_position) * 39 + (h_cnt + 39 - fish_h_position)] != 12'h352) begin
                    background = 0;
                    vga = fast[(v_cnt - fish_v_position) * 39 + (h_cnt + 39 - fish_h_position)];
                end
                else begin
                    background = 1;
                    vga = 12'h000;
                end
            end
            else begin
                background = 1;
                vga = 12'h000;
            end
        end
        else if(fish_way == 1) begin
            if(((h_cnt + 39) - fish_h_position) <= 38 && (v_cnt - fish_v_position) <= 28) begin
                if(fast[(v_cnt - fish_v_position) * 39 + (fish_h_position - h_cnt - 1)] != 12'h352) begin
                    background = 0;
                    vga = fast[(v_cnt - fish_v_position) * 39 + (fish_h_position - h_cnt - 1)];
                end
                else begin
                    background = 1;
                    vga = 12'h000;
                end
            end
            else begin
                background = 1;
                vga = 12'h000;
            end
        end
        else begin
            background = 1;
            vga = 12'h000;
        end

    end
    
endmodule

